��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�3n�� �g��簾�=8���_	rT>�n0F���_��!'�F?hq6"�����d�O,`���(�p��x7�;��a��dKm�PP�����=�X�h,��E3�������ݒ'ǅRO9�P��_͗bٖ�3o�P�Y7���k��M죘	mh����h*V(��k�c����_���܀�C��[��D,S���9��F3f^��T�=Pl40���%�K�~~!�<�Q���5FWq�9��쾙eNaaO��P:�W��]����I�s���{+�-O�X���؍����P%uA�G����Nn=d�M;�Na��OP������K	f���"7� �<���/#��`�*rV�j�bװF+~M%��`;�(1ᗠ�
k�9%#֑+y���$����0V�'�N��d�/6`>�x����r���� ��ҫ��wcH���\ʼLc%�����DO6���.0)��_Ҝ]Y����*0�o��_�B����R�94�0/�ޠ�+_�R�S��N�RH/��Ǩ�1dd�K�I�`���n��������B�a��e[��fP��$|�2�a�:>�8��s�����=�'�j��N�5@����[jx����)F5^�=��ZL�~�Q�Jj�%�9=<���:B �ؙ����)kJ�º�]�r�`�[w��,�4����"l��vW��j�<u�@-��h�U~{濡߅kxF�lS����F!�qi?	/������3�A�c��n��W�Qk�P�a5љ���kJ<T՜�����/�b�j�:���*U�Zx�n�5>X¤�XV�k���b��:0��˸1x��K�O��0�4nfb�[�_	x��O����� 	�N]�sW�B�ՇFK�����mK>�{��Sы��̣c"�Y��b�&��{��]�z���+aGyZo���-d���B㔂�s;�q��yU��B�N&5�5�h��k���=Y��"���ɤ��̷)̶$�eN�s�SSrD����D�~�x*.4��(��W����;o���ك��I��
38�|R�v��D�ٱ����i�m��='�B�ہ�$�����/���K�-ЖG����`����jt
5h�����sXY0o'��	{C��L�j�c�@W��Z��s�`JhJ�|���(ե
�G(s�$5(Dz
�[��@�7sqZDȡC����3�<�vx��k�eS���`�37�w�?'S|p�\K�t�e��O�v)h�<�t��z>_�2�G�v�/���\����?i�M�N�F���M�b,�$��3��e�w�d� �D�-R��Z8.D� ɕ�db�!GF���@C4���AH���V�-����8�>�{��8��ECv��(��}_��k4Ł�=�����\X�=�����
�� U֨����T�	�#@)�zm���W�gۊ�Q����#|Z��w4zAL��*�=9��s{�<m�1>(p��,-K�b�?�����G&\t� ���H��7��**���☿Xy���L����1�S�}�ʶ���b�t5x��(y�"I}B����ni��x����N��e)�M1�PG��az9.�^2�.�Jr�l\;����h�sr^W��.|�VbK��RY�f����R��uE��@+���͖2�?���Ws&���=���b�0*�o����npaOed��FR}�t�@E�%y:���Y�|�-�o��
�*�XD,�������R��v$�a��l�B�F��IJW����@�ȣ���
� 8��դa�����}|�!�y�R�4���n�g���sj_��>%�#0��Q2S8; ?=.W;��E�n���w^�r.α�h[�8`�F�o�1��'�hv��T�N6�-���,.Yy~E�ozB!y��LZ��iW��}���|���� p�azN��w�SV��v�eu����^�A�R�*Y�h�A'����t�OD�6���b��RGY֓��q�\��uMc���U�t2�� �,����.��1D�)��Q��(��v�8QK�բ�ɠ�rrj�5�ŔN����M�9am$0nJu�ĩ�Gew3!C���A��:���.�g�-�܀K�HoHq�(`_T�0m�I�8rn����H�0I�#���U/�z�GK�ʗIB)�W�Ų'Y�?� jr�c�n9�vs
uB ���N}N���,����۞Z$�Hг��Pb���7��*�U��1���۲e�I��:����#ʧ�����S�ME��}����Qh���DH�X%��_� ���%�8[����O=������d�l��J����o�D`��購��0R��Ɇ�++¬��h ��L&�(�˞7i������v~q�V͡��Y�U���6`�y��?����]�؟/e[ionQ��du�N����1*���OE���/�Юu�qH!(�<>�꣞?��&��r��X��-�E�)�J�0�b�iB⥘ ���C�I��j
7|�|0����mv>@�jK6*@�?�M���7r;y�u"��;9f�d���������5l̫h���9�{9�?l �9�f�Fy4�z��Zl\g���mδ{�~�����o�~��x_±����u����"0�G6��O���L�b��9	���x��kMZ��Ӛԁ�m��35ϴ��A�1%-�Cy�Zٚ4����d@�6�Ek;z�O;�.D��?L��'b��z�ݍ��8��"͞� H�}�ypZ�v޵�Zڐ�.���z�n�4�Ql�(TZ^�#�����}�$X�"�����)*��#�O<I,��L��Ex�Y��g?W����w-������V�O6����%���t�{$�
.q�6�ՠ���U�Ɩ���'������2Spv�������f��F��
�A���\A*j�y���� �c���Yщ�:S[*Y����0ao2!2CxxwHG��	X&mp��׏w���;�oT-�3����<m��?˖�9FH�-o^��r��r�e���Al���a�-���g�/�:�o�7WT_?�m !�ϱ4���|���>}̖���{*�吝c��+�tE\�q�-�!�� ՠy}s�EH��I��؂_w�!{̨�N%;g�^D�6KZ99S�r�"e:O~��� =w��ɝ׬�����gh�'"�5�������t�_{{y�T1��tJ�Vh�o>]�)C[�f��g>]g>�W8�O��j�9��T��$We1DK=�xۇQ�MڈLz�`w����ǉl�j	�ҌÿMJ0n3؈�U�i@o�&�v@?;�N��M˒��e6��?DS�U��葄�ǳg���}(�ب�GI��1�F�}���=��_�_k\�/�6�W��SANb���Q�g�%1yf��YE��mN�����ϑ�Y�㻇��cY������2���3�qp������׻�K�{m��Lf+�A�N7�[Ϯ����\���]�ܣ��7Y�Mo%*G\W	,�Fay����7�~�^)]�adTi���jWwj���1�T\���%�@��ȸ�x��!��G�l1�2S�R�`A5	��B'��_س
����K'Tpk���C�Z�z�S����ކҵz� �+gI&FMԷ&<�l��e�O�~��XKN���K�����G���=�tgĂ�^P4t�B��~:���BS�a2a8�c�oiJ,%��Yߓ_G��f���}S�۰<t>�0�o(����[M�`����1�2��(kDZ-;
J�Ҽt[щ�UֱT�zN$O��[v!띐��W��sk)���)ZaU�$I�����d�FP�a����j�%W�ɱ0y.`/�k��їk�Dhr�sa}�ފ��0�Zɩ���ͺ���ŗ�����uB�N��9%�5����|/|^4Qd�F���P�c�������p�i!)�'nffE�S�l�#'��4�s'?=PD��	_�� �F����5��n]��b�c@"'=�6��{�0{��d�hm��6IǍs�Pu;8c�`V��U�jd��.L�'���Vu�Y'JE�	>b��{�'e����9'�G�[�Vx#n����Z�S�k`��s�u\��X�<S������3��j*Y��W0��B�;�B�K��j0�<'���@ѻ&v0���/���Z�ٌ�\�2Hyc�8�S�����1S7b/�|�Su	��o]���b�~�y, }�Ue�����`B�1�x*+[��#Θ�O�=<.v��H��hQyC����&���������J�}5H�?{b�K;��T���2|�`(�5[�0����4�p�D.cV`J�"zz�*�n�7�� �O>U5�*���_	T�������d��ځ��CbC/���w_�r����?����0B�v`B�� 97�mXϞC�mf��7y��w��7u
�*��f���iu (�Y �/y�����a.��Na;T�Hr��Wָ�@����kT���}�5�T�f�7�U�����Y��yl|8YkD��I�8�"~�~__�%8�l5J��+�����pD.�BorM��I�g�:���3��:FV��������R�9���S/5�<�;t\k�NP�����[\}�0	l�]r�n���"X�O6��x7v��vq~�9�A��
 F��u<���Z�LЃ�$:���2���Ӂ�H��(�>���Ռh�C�t8e���^�u9�]@��lܫ�Qėm��$VۥA���F�نw� Ug:��x�Z>�f#=�˔��G����<��G�HP�J1������J�9�̔6&zE\8M�m�M��LC9w�]�����$�v��%XU\CH~#1�駜��R���L�!���J�S����\>j�֮�jy�;�a9}�U-���%�A��GN�a%�͞��CRn;��]^��^��]ߢ��6���4<�q�v(��d�f���f�%��^l3Z+�Q?B7?	*EO!�6���vb�&l�)�V�`,B��EmZ�Ĭo�x�􀚽С�T1����O���M��=����\ށ{�\ԙ�t.*w��w�F�!��+����qx:_o��*�R>��=��U��/�S�}t���q�b4�X�&�moT��*�{(�YQR!`���K֭[hF��7�_G�2L�^�aͱ*�e�x�y]���S/m�"C�=t��d�0�3���O���Lx�Ҽo@'ߦ^j��8��2_�1�-e`lN�����(�Q�gz�9(����;8�@���y���A��z!ѵC�G�WB�:������
t��N��Z�=>��z$��?��K&z'��U�|N��ٕN�q��6���2�:��IO�I��㛜�[��	�j`*-�p�7U�&�M'Z��p<ݫ_�/v��7���x�<��lj��i��	$���g�����C;��	��t偠C��T�'y<����l�c�r�S����P7I~��DzP#m@lW:�BkP��g���+��f�ݥ��{]#��Y��=~^*�@�-82y�z�x�,�Dr)�BR���W;e[D��#%�ɠ�М�V̢���*���2�+�3K�#Ӎ0�lZ��Q)RmeO�6����|'�M,#:č	���s4?&�Z��FO��=2z%˛\̲��ׄ���^�f���JƞF��+@\՟���� ;Џ:&������QLr��U�_C�������Y�ù�Y��V����2'��9+|����z����4�`��V��u*�&��	����_�E��C�5q�iS��Kz��!�. �5W�N6a�3.Vg�N:��2�s��/u��γ[Pԯ(} d�x���㪞�^���~,A�V�;�G%r�吊�!BѰ��ȈDAk���Ԡ!)#]i·��㖞�3X�(9-��8���nc2�/(~��[������U�I�
>%�+<.���d����x��[d��
���5�H��㚸#��V��~~:���;iT��X�Sż2��#̾����>���N�W+b�';�*0d��ֲ;��Xw�(�FfY�0,�ƻ�Zs_"�)�s�էW��g��0x5*E���\��Y*qe6�g3��gZ��D�#r�����<]�d�������I}=-Zy���$=�[S�������pŠ��$,T�ċY+3��3����GL<���z����)#4�#1��Ϟ=�%O�ǔ�}.�i7A�f�q�к�OF�'�=�C50s��
8 �NE�Ԉg��Xp����ˀu�))D�8�'�f��/0�@�U�q�n?f˴�>��4���L�(�\�TL��-v?��{J�'�uO�oQ�U�s
�mē�e�#fn);�؂K��B�q������@;���Nd�nJ�go���3�����+��o�Q�&�\1%�d;/�np"�*��v�+-rQ������u:_�W,�nS��i��E��d4����xA{\?�z#��saH>� a��H(r肧�gM;����6����	6n��ι��芺n(\�n�Ld��^]��cI
�In�5��N;�����jX"왧1I���Υd�ұ�z:㠬h8/��� �-�@B��k���R�ҷ��������0�{	GS3Ś�����ou�V�{������df��}L��%��\h"�'7�dƧr4�2�ZOji|����1c1�τ�I_��G�`q��?jgV4:���A{��n/�
%mJМ�cB}�����������L����VUH+�nwK�o�R��C�i��U��[��g����DWW�s� �_�Zn)��e��b����n��}��L,3`�40E�I�θ0"�0>�O�J�lPr��8G�q� �÷���b�p�(_�Օfw(��ج]�!k���l��D�15e����zf�n�E��Ħ��xҲ�!��j�2�D�� K�b`�����L��s�װ��KigӐ?�7Ζ}lj�<�&�c�W�6�Zv�)���`=;_�]KP���'Z �w��˒A��A3��x�"J��^JCw��V�R~�*�ߤa_T��(9^����fQA�}�9._	���j�u��?W�EFp�X�Ff����!oE��ʹ����m�a�<��0� �f�<;C��R��;p���z�R��*�h��.��� �Z�0�)M�Žc~m�/�L�_�D�N�L���p4@*1�;=�r�����?Bͪ`z�������� ����ikCp�f8[f�����p��ouCsC5��<�� lo��Aj�Bf�<M�_ة�s�}��'����w��� �fI���)�Im�c5n��EA����2HZ�"s��딢����O�ۚ��+4���ast%l�e��?8X�(���Rh��J����bxZ�w �ߠ�|���*�c��;2ʫ(�5�E��4��i�$P�Yͭ�çt�[���Ќ���HAL�r|�o+&�1S{�ERsQ�E�gۏ�# 4�n��s���_��4�%�I9͵�i��b�cg�	�8wu2R����Mm򇀥�q!��v�O�?��U许8�eV�}^`�b�7{�������C���0��vs?�����'�3��j[����[��$7��\=R�Q#hی3z�v�1����N^ހ1�@+7�)��Y�6�eΩ+��qD�M��q�cf���f��b�)�Q�kU�EA!���f�1[[Ơ8�R��g����O�[|�^X��=���g���� ]���dxp�wVdd��Fm�����>�U����^�5�Ӓ��l�4�4mM��ڷ^y���LS�B߱��z󸪕���F����O����Ϯs�S�g;5/j1���~�z`g��c� *hc���mB(i���������L4(�g�Y��1��BwB���[l����Wq8M��$ޮ��w�_g[� ���mzo�Ͽ�f�=̃��hɖ 6 �x����E��
y��i�rD�%�ҥ��*_���!j�Ɓn��.�NÓ�=*7���3k�
�%7�A��b�4xJ�0��Qgg�$9�}:�N;@�jTi<��9ǚ��w�2��^��Ԉ�G�$e��e�g�1��<�ȗ������m�:��ߊ�u$�èy��Ќj54s�i\?�#�!��"	K\��ZO��`]��G�#�?_�L���i��Y��������T"�˹�:���D�6�Tf��f����M�����J�G1^���M���<)�	RV�FYL�;�a���Z#Tw����N�����oW��.{�s�� C�N�'A��ܧ^�����/�T=CGRl�����@CP�p�__���s'��i1�%��F�+c-q��6�Jn�6��ھ�鋚���&]�b�J�d�!^ql�CY�\��Ci:��j<�2��ȵ�8޹� �87�7J��Ċ"?qr�5'~�
E	���vġZ:�~��zC�TvJ�j�e�c�0%�ZO�����h[�5�U~++x�*B���Q�&��4��4�&�e��B&�n`=�e�(��Y=���-S����b64
Z��3	�����'I༥���pߝ��<	���e�FJ�nl2_��$p���b���w(�Z�`��D����{T�x��aH�6BXI��6�b���7���&bƟxii�ԋ�t��i@1�hr"�
��~�#���F�����-*!ӏ.�x��c���5}$���M�ᢲN�>�RM�:������h�	�j��3��""06]�c��!�h��<dR���$Nv�֚��i�Kj}� R�r�q��U���\F����OR�m�ܧyƃ}+h��ְ�K����$�I6�@�q�j������6xT|����N�x*���v:�uu��f�d�]{�@e�=�����]����7��}r��g{\���{[��T��˱���%!o����Z4�qݩ���7~��(=�v6�j�4�홁vB֤UK�"����Σ��&!��� !|�[��tP�����b�7ן_*�[�^��AP�B�oy�b9!ɾ�>����T�c�wO�f�G�(q� A��T?	NH���@��ҧw?���A��"u���:�b>��UŏUE�A�� �b�bRd�>j��<��'&^�ǪvE$���/0�*R��z�*4dh���D��(�rXq�� ����]�h�~9H����^� r,L��j�J7~�b��~��W�=�ha�� ���
�9aK�;F��S�4�H���PpbmN�2�F3�JyHPM�P"I�{��E0yo�Ӌ ��ehWߠ���3_�����OȆ�f/��PY0��k�L*M�A�@�.>m��L�rW��L�'׿�/