��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�M��8Wu��_���"���8;�Τ� ��֑��I.5�D��{��	˚k����}Ҍ}F��n	�׷BX�P�;B�b��'��H�iv�Y&����j3X����-�����W��;ح��@�Wk����*��0� s�����شC��0�P��q����������J6�v�׫�q!��������>��!"Do�Q���,g[���a!Qt���c�)ؑޤm��r��л�Hz�b6�qv�������M��ŝ�9�K7�;��鮨$�X8���c-�E�h+160��~%�^�Q}����Ј-�CT-�Y�ՙ�V�o�e���ހa9���D������C�Un���ګ��z�`�����(QW��h�d<g*N��q�YH�Tw�ue�h��LF�+��*�I|$.�J��K�5���v�9��������6.7����LH�椓��k6�F�C?�'9 �0�(q�^`~Qux�A�K���@`���(�VaW-�$e����얧�Ƒ��$f�z�CO:vP�4_����o�yU��Zw�Xj���O�T/��0�c<�4&��3��#�Vy+�+�yU-k�OP��Ρ�DÆ���s�Ԗy.1� �ʄ���Ύ[ElS!�(���H��W��di�Q��E�AS/N9�l��L�w�b��J�::�]~�-�f�P��0�X��B�㧚�>��u�����w]�r]߇ۅ|Ie��%�u���P�*{�se ��!;�^5�[�ٺ�Q$�R�nE�F��1A�x��kN����#���lv��4�oٝL/WA\���Ԙ��k��[�E՘��@g��9��<�RI��Y�L{ʦ{�H �"S�g9�2=M����]-N�d��.g��{�!�%�l) X�|�4�
�A��&A_��u�b�
�
=�x=�0��"��P���F�H��ȍ栄o����F��h��dʝ-7��z�3�-0e��`>E���t~��iu������ğMF�l���@�)�wHІ�˰��ݢP��h�3S�&�h��L
b�u��%�S̴W�82H05s7���{Ժ������w�ɨ3������.�p�m�;��c�G^M���(f�#��I�/�Q��g�s�bs�v��8_ʰ����3�z=��M��p�Mk�����G��\��-o,U2�e\A��:~ˤ%<��@z$�#k)ъF;�Vj���bV�*��t�1Fa�����z��T!<��d+'�Aq��pJ���9��э:���s��F�g��)�������}���qW�haΖ]*C3$�&����^�qx#��6PK��j�	�oo�*)�E��hE��>�lVp�\�<�NCr5��٠<ڬu��V0�3�M�.d'x)P`�D�cu%j�-W
T������'`:��A`��x�dq���LGN-�3ͷ�D'є��A�c�V��@a��`Fl�U"�?�*E��-riF�ʚ5)XߪO�B L�z���Ȑ�-��)�A4K���w�l.��(�Gu?n���R G��0���q 9����3��~�W��红���T�F׎�O��o��::D����n�T�!��8\�X?����7���� �b:�=����O�)�ޣ�I6���I���`8�";>��f�ٸ�M�q�
��]��t��6<ח��_�ƴa�e��p���q���.��vF'plR��]B�r�h:��ﴷTt���4�[G&3N���C@ O�V=�TI��V`V�k8��]��M:���~��ש��O��Ӗ@���n��h�/T��L�N�4i�x�Iv|�A����̖^~�k����c�@lW��	Q��.G�"C�e�b���5E���~�%��i�@�]�ӽ��ր�e�&���\� �{"R�@thTC31�%(J���������'滙��Wb��Ł֫�2�?�E$���!B��s��o�!"|]	�-�G���T��:e#�f�4cK49���v�B�S}�{�΄����r�5���<��-+����4߇�r?o	넆�L,��:���-��/��|8��cP��}�I�A֡#E��ȼ��]���L���e.�O����
j���}QH�-���N��M��U��+<DT}c~����'4�Q��J��lZ�Bp'��#g$�~�}��yAI3�T�D:�����4@JRF�"`a�M<�=��j�y����(��P,���)�
���+*�J��	c���fXT�����Y��)���A�E��NC߹���b*�U,F��4��D��r�O.�W��]��g2�;��];��_���i�c�&Q&Ee�f�O�6���B�B�6۪�ۺ��a��s��	��T&O�z����¼ =S����y^:ᔮ��Xc ;ɋ5r�_*�c�N!��Ӷ��^����v~�1�w7�`Tm��j��nȾTՏ�K��G֒ɪ�@��o��L��{��;�4�,lC:�
.�Qj�xg�28��#�:C>����oQ�
07Sw)�nF�x2:9L�뻏'2E�>�Ұf��trJ\�OvA�iM��F���B�����O5z�f�-E���,��t��7��s[<J�������\���e��F��Sϑςƞ�9B���`]��+M��q�m��$V`F�0#\�~~}���\ؙ���'ђ�ߎ�$Jˇ���c�����\�&�Mj�~�n;o!���(��u�_/�X�jw�@06B/<��g��-2eE�
���N+ep!��i�����=����8��|�� �jȹ�-Q����]�v �)��NjkLV�e'�Bo�=.Q.t�Bw*��&E��b9���P��X�I��}V$�Þ۟������>J��� O|���2/|j31�Uz�Si���h�8�}�S� e,|���$�k���O<�͛`m32:n䂙�������F��s�Q����pu㤿��Nԛ�<�1]sa�9 *IMf�.�W����m�ܾ"m��G���j�z�Y�=:�9�(�$.��4N��r�nq�I�*{[Ka7��?��dK֯IX��w63�p�i2V!!T�jFy	EJ[*�(�v�Gdޔ� ��`�!�:R��[�~+$��'ah�ZU8�f���k�����ĻK���w�0·*ŵ0�r�eD0y��d)[1�r���
Km=��Ƞ�o�x�MP�����1Q�z��9�6�������x�U��+�
(P�����������ԡz�š
�+�D��s�CXx���9��T}�~�k*/7���@���m*U�42oS�.��E�RԲ��*��Ҷ�$��m�}�+�Y����ŧ$�I~)(�����*���=�C/~�����z�v��Erq���4R,�R��g7��U���o>���9a�f,k���c�W>�s�&uW�t�;�,��?�