��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ���v��+޷,'����]��<�GN�J���Enx�[î�yf���W�?�#5H�#���M0�����Z�����T'�Ȕ/�ϵo�;��T'-�}W+�ա��U�5ٍ֦}�O��C6�xp���ة�Q��)%ku`9t�֨�68����%��՜+��WO�`�UֵN=��o������f���f�Wc�)�y(�{�qt��J�6b��Bh"w�T�5��3�{��*�C�Q��;G�b�uY����:Sۼv�,�%������h��D<A8ػh�}�m��ҝp-�A�U<�7��Ec���i�R?9�6���b���"���s(�7o������޾c�W�c�Mb>'B��U�;�����5��O�!�.a�;��:k�5>�*��q]	�l��T�ʚ�~�z|p*y��Ɯ/�YIP
�F�1�M��Qlօ"5YGc�L�ړ���v��W� �[ϝ=��f�i�b-!F�X
C�e�R��֝ȭy���~�C,-��F�����l�jk�����ce~�m����bG6��GO��V6�0��<�:}���"��?TM7[�r�� 5�Ovf"!�8N����"�2z �'XvqG�[�o��4�X���ԩL��i�Hx,;���+�����}i��Vs�A�T��}�b�p��n�b5�� ^��8kJ6�Ʀ!���'�Fr�ѡ��	zih�}׮L徳�!4���8��u���j����^t�)L����]��Һ8T�m�z�p���BSoc??��Z�"sv��T���-N��-$�"O�`0$
��P[�b
�W���m�'�Z��x!h�;� 9ج蛫���r0kC����	�ˊN)<�~�7~/Q�
�d'��]�y16`҉q�O�U<�Q
S�LZf���5VE#���<�������΢��%���a\F>|@�#��gGA@94̥k9v1чT��e3$i��Y"�_�kM��CI'�x��32��j[�	�U 
/���'0h��/=��!X\td]�#��b` �O4�+-����s7ݒ�U��E�>b���Zu�^�t��=-�$H�ԯ���G�2x)2�4�:�e���̝d�Y���
f��c�K��5���Vsy��Vd����X���8��Y�3��:g�K)ۻ%Chi@�����:�A	����Ba܈�EO5\���<�Ц�F��S.�w�M�?X�J��t�����Z�Ϣ�87�F#^�_�J�s����1t{S<,��� @3l�T��wx��Vp��˸y��Ѩ<��ݹʼ[�4���Ti3����r�J�ӕ�Xů_ -t��)�A�Z�(K�yC��v�m��������5&8Wz�����t���s��׭��T���?_�(��@����i�b/���j����VW�1�e*�Hp!���eІ���ֈ�(����S�^�Ow�,����+)�{d|vz�F8zm�
���(W��+0��s�W���5wK�s�&LA�����P�4W��[�]��z���/�&�1���d����Ŭ'r�?����YAy�X��\�%+� 9���]����a
jXEs�F�5e��	k���#|K~(���&���q�����`��:����2*�	�o�46��(��@� ��.8;s��e^>M.�������X��Yy.�vk���)��� �Q��JH�r��(7
�[܍S��YqlzEw_U?�^�t�7V\��(���f��8����2�h"s��@ET<����}�"�]��R�\b��4tΩIV�G\���R��tV5GC����W�p������PxR�xW�H�p��) �m@�C�̀ oEel~�����0�w���D�A�������qg�<�{���:�	�S:q��?����6\�y�ߩ0�Z>*����Ļ�I��{a͆ߛa� ��c}�v��Lˋ3����H���#���c�#���Ԡ��lY7�^�\���cgp(yET�+Zx�}V�T��V�z�B8��V	�@vq��7��5�M��T����IW$�L��60q	0��9�-���JNaF�/�ms������Y��U�����,���9b��} �<,��q������M���̛X�J���Y���G{�(I�C�|��X��db��T��摸!WMA����ŗ�N�v:o���;ߗ���- ��שׁ��)Wx\��^��5?yj�
7K�V��2��X��P! D��J-�Ro�y�<$V��7.V��� UX��$n��2��+�� -^}0&=\֘2�A�����*�ϼ�P�$�`�#f��>�$��v��*�$ܙ@�Ŷ� ���D��b3CR!(�����_�JS� /�	���G�iY�`��NxZ5D`�r1ӪN�B�{LlX��Zrdi0S<F�2i����q21� �#]av��ܵ�A3���
��z濟�Z���� v�y�^_翦s�9�Y����kA?i2�	��s&jûgT
���W�ޅk�i�����G����K������7B02���D��n�IZ� ��wH��lR��M`�4�����>t1��dX�<�#�o�A�����T0?i,E�yŶ+޲�|^M���~|�\��/�{C,͢k�z���mN*f�PF) msx����[���]{J9�lU}��$�� �i�	��r�S7xh�T���FаY�Q�Up
����Q+s�>-C �9A)�n�`4�W���1-�tV��\]�-7�ȭ���\��S-��k�ǔ쨎>��۽�����m�Aj�;�� z]�g�~��(m�u�U���Б/G)���Ŭ(P-��U�wÜ��jw��G����S�i���ʨ�����{�b;9�x}'K�m��$z#�-��Үd%�(w�O�)��\3�0i����`Z���}��~	�!�Lѫ�x@�.+���LSٟ.+k��E��-L}bB�E5��(�#