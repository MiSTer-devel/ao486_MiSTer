��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��ՉN�*�s�/O\4��>�� ��6.iT�<�����t���K�6���NԲ��/�;��F�U�*�!���G�@}����M�c0�y+Gp��!��Mb[�>k��,�%g0��\�,�󌱭z��	_<-"��A��m��	_a��,�e����/�x6$N��H�T����aP8A��,�<jbܖ>0�ܸ�-�����I]�u7��-�Z����R����S-��ۈ/���U�]��;s� ���B]Bi�@�wZ Ȧ,���{Ȫ	D���'}��2tU���!�C����!�Ң�l��/����=�u&d;�`_A)��H 9�h�U���-�y>�#Rn[����>n�i��i�Q���$�}GtT�h(>��`�����,�1���븤Y�R�h�Le���hs�����C�w3�Ʒ�?o��p��W۔�H���T�w�����T����p1������ �h�5����"Y�x��̪�y� 6�u"��l�l�J����H�K��D�E�����&�u�P.VU$���p�L�N��iY�'d�q�Y%����7V�e���W�r4�_�G�F��
$ ��Ϛ���GLs��ZJ��'�t?��2����*���"��ق<���N�Ai3"ﮏ�u hh�p�dC(�Ƕ��,�9�@>0סDM����_N�RYE9�P�ڻ�,Pv-�fe��F��k��pݪw:�Zԙ�T^(P���R 1ڪI� ���jC9�!U�����d���L�)Gh�#;�-���[��ϊ�/p��ߌ:y�1@@��.�s��a�S�;��)���t���M�!n �