��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�����`ط5~Yd��d��q�F����8M5'�d�la^M\q+�s���EB��F�mR�[����V#/�.@��n��&6蒸r��M_�?�-.����#�+?��i���҂�_}�N+�9� %�z�Q}"}�=vF~�QO��ʛ�V!�gI��g�b���E��7G�ˠUe����$�\���Ö�:6�1OdPjmQa����|�o_C���=�-��`��qr�z�����Fj�*��`��C��@�Q��R΂Rm�߁����Ke&I��p��/sQ�t�fsh��y]]�(5沰ׅZwk��m<W��w�:\��PA�<�#�Au����Y���N�AƷ{~�����"��e��a,\�CW*�K����W��b��'iSo���:��4<���,���C	���*���6CjJ��Z�l�=�Xi�'���|`�H-4
�7;G����yx�M�0$-����sv}��k� ��{�D ��B���̥�x���P#U�������<�u���G�
$�����=z�����7P�e���1DYn+��pT^�pK����4���q7>�5_1�Ʋ�c�a�T�K.Ą5s�����J?6�-^�7Ї����WF�G2���9���}yw��eС���A^��%�|������џ��(��~U�(���JQ|�o�>�P-a�3c����g�����������d�ˮ-��A�ij�'�vI���\����`�8u�kT��F��+pQ1��3M������B�ӹ���Ɋ�.WN���2S`*�UI�}�p�}�($�*c��7�Zr%E�[��#)���1)�  �u$n��I�0�� ��%�E�L몧��y	$�ܧ����!��^��%kӠF���GwN�H��y��e'Ų����Rq Ɵ%Ld��x�fs�x$aDK>W��m=R�<�F��,E�<l��B����j|�1N��;7]s,����6Y9��L!����/�M�ה�2a�����7V�J�A�vcL��N�L�������*�����},� k������;*oe���}��8ȣ}垜��L	�+EԢ�<�ܻ�Q�Lt��e��f��Ɗ6D���=]�L:���XPMf�6�is�z��b�st��
^k�P�J=/L�uO����O�'��VO&�Z�M�ʤ""���� ����٪H)%��d.0~�9yo��]�x�۾E�����X��IF�Oش�<:�+�4*x�r�O:�����r����
���A�x����N&�I��gʁ��H�9)�6|�5{��P��B���{��������L��m�O�T�6V�{G�������^���B����u�� 1k]���Gw�#�U&��f�gS1���c�	%��s\�i/_P0伣4��c��.|&<bŬCmJ��'R��7^�bM$�K;{����M��8������!�=Q������#iSi�qq}�6z�R|�{IH��+��_������92M�"'u40A�ТA��� �wP�	���T���_�T��F���v�ӻ֭�I��->���"�s&
���%����5s�Zz���b8��г<�����[LA#��ä%�q��|KN]�7X�� ~�0�<�������B^d@��Au�y���x����-�P7���]
�b�2=|*���Y�F��Xؤ��Y��7<9����7�#���l�U��� ���a����ȖyLڣ�jR�T�yز���q�rc�04Y+q���2mm,�j�w�Ӝ��1l��|eY���y���:n�Kc���-˳@�'U��M�5�H�*M�����  ۷�Sb4�~��o��c����T��L\2#t�5�A�gP��]�?�p# ����X�9y�!QC�[�s��\1�P0�?ev��\/Ǯ�q��!�M΁݆������䋡扩�WϺ��ͭh�/�P��g`
*��zI�8H���7כO*��0�X6D�ڶ�c.���' �^�l6���	����+��� �M��x)�|�E���&N��m1�`�ݻ%y0�,A���_S�ZM���6)��7����\��\Wf5Z�-R����"���/}��ܫc�V?"JWļ������+��VW���!�a,-3&7���+c��f���\8��<fR�ǐ���B���"� ?y������ ���A�Yߣ=�}D���|���,`_�H�������aw�|-$x>�)'��)��X�F P�v`%����A��(��Z��%��U+JZH~X	Y�w�`���H�kӅh����j8�(.�ă%]Awg��t���ߚ�h�� ���?(5�Py$��"h1�[(f�R��F5؜�}u���3�t�X�M��З���f����g���+{|��,�l�djwAц�:�Z���:}����وz|v�b�nZ?.n��@��i�2�0�=I	�� t]�C/���C3/�h~oav�J�j% �J�,�@A!����|�=�s�-Dd����ע�#\n�N	�z=��yZ�R��B��J+[��ؗ����8'nt�5��Q��S�h��2��N��*plT��R@�3�9�p�>���ޤ��H�H�~�l��N��t�7�~X0Q�N���\�i���4�=f�L61���V���P[�L��&��  T�mOTכ_����Y@���P�����y�?���U�����Pt�3;�3#ru�&��e�Z~�]�<g�(��C�aa"����-C2�^|Nsz�I3�O��"%�..[agr��$8��<G��U��ӎ�M�I�Ώ*2����ȫi�Џ=��~�"���$�1!]����������[`�~���h�2Ф-��S���Pb o� i5m��X�t�I�x��c���lu��x+�Ak傢���K>���5��^!Lu���4{ ��ܳ�O��3w����xnL��KY� ��Ҿ.[�����$�n�7D��eE�{p8��oU_~�W�	��3�RRkT�6�7�x��a^��A��P%w��	e�ϋ��9u'.�)�&��ئ��;��k��z���c�{�c�^�n��^�J�Ȏ�_��_���{�s�>������<?Q��*�A/��<��G��
� ]��C����G}��?�(�lw�T���caOmY���󠵢̣-�1ߢV#|�:Ԗ��Y���Xz+Bi��<cg�2ʴԟOҁ�5���;:u�`Ffa����;9�� �tLuE��6�����%�=����Eo"�ܰp0���q#o qa_�WI�+p5U��ER��S|5�f��J���A�v�U_.*m	�a�z�	��#�K��N�s�ߧ����S��Dz�fX�����M3�=}1�(iUG�.2!��@�y���v�������Vr!�GJ�5r�`�6A��\���Ħ��^�A݉���3n%�m��7���
�x���8k���fDrm�4�l�M_=K=��n6���W#ྱ�6�� ��P\�L�]��ʂ�N�|�`��w�T��#c���g�̹�O�6�8ON�ƀ͟��֘�)��d-b�T}�d���hq�RZ6��c�ǜ_
���3�(x��OR����VK������&���> ��$DNU������ѡyg�م�����t9d=� r}�lk���S�%xYY�zz�o�4K}�蚂����h�Xŗ�|6g|曑�ȶ�䊬�s��_iHr#�S����h�f7���E�0�Tm>�o�Mռ-͐�����b���1/r�En� ��CM_�h|�
�vTv�_�x��]C��<0d�ኖ�5T��'[F2��k%A]_���bۜ�m�0��S��|�C	p��v΅E7,��.�dh_Q�����ȃv)�쒇���3s�p �#�@�gZ�g��R�#�9ձ�"�U]�g�=
hkwj��
��lfk0yH����:��W
'����	6������a�2
NhI�~d��S�T
��h�߹��8�Q(�#�N���.��=�,ea���|yl�3h&�����JH�)ۉ��Ӛ�ݔ|tH�$��*ݛz�n[B���T��np�(���b�����|��m�"��������Z:v���'.P�T�c��|��eں�P|�����81����'���g��=��0��o\C�Ы�#�Z���(�Zj2�C|�nq������C�{'�{|[�u��%���N���ޤ(2b��:��g~6���ݖi��n�㊸}�<�`��D��X�[��Q�(N2�?]H"�N"��lQ9Q:���C<`�e��g/��=�KG��kG��z���S�c����ňjR���������+��a�O?�����1�ث�ae0�x �u��3s��A�3,�~KG�L%ecpI�K�U�V#�$�֘��%Q�t�������`D�o���жuiO0�jQ��mƯa��V��K�������eK�Wz=��6�d^Y�st����Mњ�t����}�}#�ٚz�,'�r���h�^�}����r�?C�_���f��O�{˂��c��ç�H<��=�WRz��`����� 4�7,̬.�� �r�� y| �FY���箹��}�IM�Ԣ���)��Aq���PVn4(��R��aj����?�l9���g,A�텡�~�Hg��h�9���z?�f��{�.(��JG���
�O%�׍�~���2��*o���s������)z�'dV������z�wx�E�RP��z�4�zB{��B?�}�����`��Xן���	ĩ@m�|��S��r��j���ҏ�f��.eN"��B��]��E���d��{����Y�F�!���`s���Ɣ����0��j��H��pY-Xi���h6q����|όsE����P�֐]�,�{ܦ�'Ag2�m�I