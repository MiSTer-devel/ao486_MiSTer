��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ� t���=?�'���]���y������/��? f�'p��O���=�z�5w$�����=V����Ӣ�.ny���Β@`&|����]'/�._��2"{����x��&˯�����5r�<��_S���0���4X!����^a4V?��>�����h0Ĺ f�$h@s�}�q�)�1T���hK���앹D��V�:�� SW�:��!��**�֡oe�!	|,�k��=�ˊ��o�P?�2��y����������J\Ra<�#"o߳Y|�u� ΋
�3�O-�`���$�D�����y��9���օ��X�ϲ��RH�yE��> iI��Ii�vܚr�~��	�%��������#�D�ω#�oa{�P8f�����QI��g�#���]��"59bnj�Y�s��3(&�P�j��j�f����h�,!:t!�*� �9��:���rQ�<k�[�P�A�QZ$WZ�緎śWn���Y8��!KH�p,��U�'�߲�*I��폌��o^��୹WeW�,}|F�p��^ (07�&�o|q[�
0:Ӳ��S��&��h���t^���OC�.����+@���S�ǯ�����#�g9�dXpd��vGS�v{h$� �SӍg��o�X=��I`��\<DH���G��đ��c6��/�8�	8PDɱ��[7M����` VO>2�;���#i���Xc��H�T�;G�Jnn7.D�;j4yU
5�O�A�s�� �	���%�� �/�m ��*�ݓ�*Lc��,���pϰV�=O��	K픜F�L������i����bU ����p��L��"Y����*�� 9�JF�İ��om����9b���T����7��_&�H{V��e���6�[�I����i<0D[���Q��E���e��[�^�����ɲLns�<!��@������V�2��9$��m�l<|<]��Ј�Z
�5}�_�Q%�^D������_���-����ˣ�G_ƝP��DQh�x��oV��P�D����t,~��o�9߽,����tD�,�G	��5F�f��B�5��U	�:��U;���Н�r�}Z���.��Lr��Pޙ=�:��$�R�f���e�aa@�Q�I�t9b�M��2��A8��h���8�~�dkp�fm��bE����;V�"!�cW�a��u��@�'��U���$R;]��oܘO� }M�ld6�	��Ӱ{,�w_U�����f�����r�Q�ߊ�@������� ��|'��U�Js���/�WM�l�̬6~I@S�#�^4���o���ޱ�זtN%L�iD��A�n�+��N���j������ ���"��nL��i|�/"�]�����~4}�2��o�N�[	����L���j���S�NH�*��X��kZ.��9�i�	�S�fg��M`�{�[���B.Yj�)�������|-�������얭T�ۊ�Dd<4U��mŶ�[�/C�C�9�^XH�YV���]����%����Z��z'Q��+���mUN���*%c����0��$���7t���z����"~d�Ro�z��@�Ks9�ɶ�3f�O��5�2� p�
�X-v��/o�n�Д�,�0��$�t�YP�)_w�Õ$^�d�|!_u���5� ���"�b�6�T�D�%'O`�W�?]��m*��	{��&J�
�f��<�y��}�k�iv��m�(�:���9����[B�u�G($/�=ah}I����9[��^��>|,a����f�\3^t���a���*JQj���߃ _�˛�w�M���.�L�)������1���u�Qw�E�a�lp�E!O��}2�ەp���yN��V�B �^Uf>�Ԓ[OmA�^6z[mJ0�Nu�LW<�<����Z�&�N�7��c�3�>Z`����D7sT�yx���J�="��5XO�6�t�aK���HQp����4����ޅ#ztU�}�VK�/�ks��DbP���0mo�.���0-�-�FZ<W�&D�E�PVL��6�^�n���(��ۘq�-���`ǡZh>O�_�13î7.8��鄍�� �;x��\#*�#U������n?:�T��|��a��N�3�:T���r}.�f�L&#�����S��r�~ �"��oe��^�xg�y(J���~7�+ �
}�EjH�)f�"�LIǶ�e��ul��Td~�->I|D^���A�Z��� �x��]?�}��������$��Y�/Z�K���ޑ�^�ˌ�����<��d-V��Z> ��R�=�< ��-z��/AB(L��O`(*�ZA�Q����'k��yDn��v��\f�f�K���>�t�X�m�d�^������t>�M}Ȝ��e�Uqv5H�2��-�k�_��Y����\��Һ[iu�{�'��o��Qr�1ӫxЉ%]����j�iP�c0����y�tTq��sWL�g?�5dҤ]��{�*y6K"������eSWs��r�2qSr���#��C��SN���5
����6&#[���K�&�+��$�/�)Z\k���U��K@�E!@��>?I�S����h�=�y��r�Zm�vV�@R�3c�a�%z�9��XU'&V�8Bi!�Qy�����zV��c���:G?�����d8)����e�ڥo�p���)	4�BZ�\%J��5e�y������\D�*թj>�v˅���A�xӇ77r�k��2��0@Bpܱ��������;� *�oOw-�X!-~����v:�q��m�8bΜA�D�,8R�99qR,�;���l}�5� ���Ϫ 6��{����0��Q"��2	�@�����Y7e�+|�T����ʮ�2ؾ/m�\K��4�]R�����O9)7$m`	e�;�<��ۑ��5�|B�
l�`KW3=��,g�Y�^ѕ<����'�׀���B�7F>J._���yO,���������|f�1�wx6;?k2�Q���9����̍o�ѿmR�%�Rz���k�Cb�L�'e:|W�u¿�oL��7A!�EÃg�������W�}W���7��>4QӒ��m�oi @��\�dtmR�V���"'��U��Y��EwS]l�ڪT��t�he���E��Hcz��n׿3�G�GD��~��NAn`uS^2� U͕�wtXg�\��ʜ!4�@�|�$��d�e��U�	g���ES-�BT߃�2���^
F�n�Ak,tއ�8�D٥�!:=,�A����D�������D����W�';�lsM����Zi�+��������ѐ��ޕ�뱾�����2�5�o=|��F¢t��M���έ�`���<4����D�f��k2r��m�M-�|��-��A�I$?'��5����s��Y|U��Z�$OyC�`B+;���3䜂��OG�u��	δ'����c���1(�����)(0�+��.�owQ��'p*xL!4y��0<Be̡�K�Nd����0��9�eq���1��M�3L���3�
2�Y���8V��;E�/Y=���6l�Vl{I�}:�^)O�"\��3,-T71��xx7�~Ͼ�Qr��#ZjW]\֫�B�V/f��17�B�og$�d���f��ɻ��%���؅���6���)�_���8����ڸ�<5y�[�X��ƈN�U>?yf.��H��ْ��(��O#�?��[Q�f�N-
���"I7�"�&�2I�݆�v��s�դ{]
ՃhZ��ڗ4YT���im+��8aK~��x�c!Zއ��ft��A\��=��w+>/!>�$�I���� �=E9�ݶA�5����Q�Z%褥/{"�N9-;�Yّn�b��K-Q#��&o�B�R~����?6z�c";��BA����nc`���l�tPB_6��P��8L���Zԫ�'�xG��/u��^���M���
�U��)����g�K�:(��T�x�o�H����>Ʌ�ZT�W\A������蘗��#�
�%Q/���y܅�5rS!��[�>3���J�u��_�y&dyDm�@;�0�������B��\������
�e}%#���a?�k��2��V�WMuƳ:�Y������������v%��z�/F �O(��Áu̲�)7�H�]�7��#%`r�{���:�����oh\>���=��Yլ���F7�!�-c>K���Gpi[b�x�&���q�պ�5n(^�e��b<c�z�Mm�p�"e��vy�`�?4���8�,uJ����7���%�N��{��,>���W��l��hu. �==P�Wa�<y�eEc��g����͉ ��Ɂv�ò/ǅ��:��Ø�S��5v Ue�&�_�U�3W�>���F�P�yͫSF 5ob ��B>8h���������{�XH�����Hb�{��~��E߹SЅ�r���}6�$���})����G#B� �w�@����AU��l��d����jV��{^�:�����K/��1����M��Z}���2�����;�f"wS8����=� u�Un'm�*汑 ��61A����ƃK�_�B��
e:w7��gf��ň�SB��c�t =�{�c�e�5.6<�o�+�g��кx��t#*L�@3*�o�-��́�>�`�| ٵ���J{�ݻ�dY6��iY���4�
;X���h�^W�/����Ϥ7f�0]#xƫ����r�~�+B�<P����Y*Y��QDѻ���'�w$]TG�P��< ���i��:$�&u-�Y���ͳa���B@����'��V�x~&��Ç�칳v)�z�Ɖ�f�Cq�肼��$��rM$
H������Y�	�e����䉡b.��^}%�9�ƌMH�v=�l=��(=�DN]�CeF�M18�?�*�yz��X���vl�6Q�{�m��v~s�'^*�5A+�g���ً�n�]CZ� �����H!E�b��@��z�{"0o-c��*"�*�qG�5��Fq�{�)�
x*��~g��q��Ut�Z_]������Ǵ4�cm��l)��[ѻ�Q�&��31ezf*U�F�2�R�^uDfG���O�����"~�H���y_gK���wJe�x\��ꪢBp��̎�xQ$e�Ֆ�[��vXM:â�Ier���g٣Z_�t7�j��&s���[F����p努�C̛�7Hٴ�G�54?�X�{nwbȳ=UET�R�'�3{�)CL��#��lՕ��{V/��r�a{��}a��͆/
=?9�A�T��@�f�:u6���>*z�|C�b"����E���x��ME
5�,�x{/��L�HTW� ᢨ�E��[;Gœ�B�ǟ3�B�Ǿ�҉���4���\j?�y9��ɨ�����؆����0W��:������|�m�*ƚ���#�]�Q
���G�^��LY`��_��a��ɛ?`d��A���F�}�e�>�qu�{��tq��p��iF�ǝu���Y*S��]ɟx�x����&#,�ˬeP:b�W�h�[;���.<);�b�2 8Ew��w+����wJ�F��ePD_���e��/�>WD�F���q��9��x�ɝ��qhY�S���(���Rl��g~c���V��;4���]޺+0�i���9Z�Jz�ņ��˙r#���� � �4��!1�L]�:I�5X=�bmK�M��RK2v�������u��6zᴢ�G�r.4��nbU�M���s�6�l�yx�n¸c���h}6�O�
����fo��#�g�s!f�L	�������~���	����/�U��~��.��y$s ��f�$���F���V�*�����t��Y5����5�C��&-V�'���?	��%;u�Y�Ol6��K�����sГ��mu�82���q��,P+O��r�c-�\����|���E
���& (XxU��B��r��hK�@�t�_6���QY�~Ǹ�������������RAh`���-�����\��#}Aq��!t�l�\V�sk��\	�+�B��Ky���=1�
d��B N׿%��� <)8�7#G�V21�ʎO�s�d���9_,�������Y��x���}�'�T���3c�6%�<R�"
��H^���f�Dn	�Oy��'KK�qc1!�×����'��� ������A3a��(�??Ý;f֦*Dk�;74Jܴ��f�;2ߔ?���b��=��m�ta�����=�C�3���/��	���T�4�[ͦ^�Ac�K�LSf��l�8KB,���>X��G!�6�dB�+'Ew��IO������Z���`Y����(��
�˿}6i+�%�����b)ᠭ�����|��ݑ^��+�B��g�����4/��w����ŋ�� ������b���,G^0�a׻]��	R�`�lO�	y��P\qʍ��:��O��]A���%��ݬ�f����m�Ny�5����@�}o0���]���3���ζ��]�	a�m�7h`/B]�X%$i�C42��?���l蚖1��,�	�g㍛�/�R�,��`�*�v$u\�Xy�g�s�؁vn�BeF����'�4ګ�y�'"6�)7�&/�w��QR᧕����q��7ݴ�O��3/P*v{�s������f1,������������gje����Y���p0Z4!����@`���}=�{BFF�����i:��B[D���,���$�s@i��C/9�OE���S�Ÿj�$t�?I�}83y|t<i�y�l�U�ڡ\�W@s� ��ew�d�愣6B� �r��q�	������`wϙ�Eg��=��`vP��=E�����������>�t7�.N^Cx�����[��>�U`6{G߬?2Ɔq��'"@�:�ʂ� b�3��{Kԕ����J�O5��M�T�ÞvHvit��iFR��!X-�"`�����@���Fjy��
YѨO��a���<r���;tk-�O���wR��4£�z�����K���k���@��#���:������~���T���RN� ���2o�Uc�b���ó/-H�ђ�Ӷ����T)�w��;�)�͉zҘW(� �0M����pG0#�A���A�'�?bs�������Pr��=�O�q�Rd��ǰ�>sֿ����d��˝�U&\<s�ԩ�L٘B~�T�Fc&BN���^��n/�6^M6_*��J��$���,�^�z&�j�
�g���ۂ���W"�bu�~ ���W?$�D��\#��w��-F`F�%�X��96��E��LB;E����L�,SEw�s���w�l[g�:��<4gm3o#=U;7����|���dӥVs�G�d	J�7���w�/�D�67�X��f-�QU���rMtmfw�HP�~1�J��/��S'���)l�B�ӟ	;f����qbR<}Y��N]0�R����Î�a���'c?�e�t�k�q��Pm#�b~�"�D3KLW����Һ�ꗍ)�mK2�k\�)�l1\��ߘ\�g癫n��))y��r�i��K6�{rC�3DF~��<��`���'��Oe�Wf�dI�����WMY 2��U�9G�M$�����xI����8v����|Co���]�gT�\4�M��|q���F�.'��F^�D�d����/R�h\VK���>A����*���A�s�Quǫ���2�}^�0�T�B�U�PBp�t�v#6v?��A���S���1���BS�N��*BHY�Iy���>T5�F� ;����Eҹ�lu��]�lpb�G�A ��S�\[����\��dտ*̙��޴�����K}�7����~���ぼ�b����w��y��:�W���W��%��U.+�}�І��V��>���r���N�4�v!�W�}������Nxe�xQMSdd��9eK�<�����֪R*��7��c��/�l�-�f:��Ͱ#��T���mY�_J�*^
���S�[���W�b�c�k
$c	������������x�]E��"b��d*$��e�	s��@�W��+�1��9�2h���n�.��(�ڥ��HOJ3������b,Y�A��cU;9kh��@Ѻq��eJM}�㥮3���h��Z��aZ���m�t6���­����f��Hd徦�D�i/�-9U��5t�c�&���/�3d�M�o��,X޿̝�n\74�,U���j>�_M���r/��qҎ��b�&��4Ķ3#���A:�Z��'bMo1���%����i�e��gN���~:T�ū����	��g�F���Օ��ZX��]�0�`�$���]c�{�)���N��0A�u�˗�#�Z���Ճ�c7���ސD��9T�Z���g�/��w1�(E�3ɡVu����ZO߿��d����8�ƴ�,Y:^�Z�^Z����Q�����=IkW�%�� �{�j$v��)����&��a�����O�EW,��#�R'�OdZf3DT�Hck��HH�8�%����.�̿;�7�W�F�	ڝ�h�0h��_�s����#��m����\\���h�~�����"��}a��>g@PB�q�2
���>�N'��`��������6:˞�g~N+�c�=F�b]_���#' �͕}W3�j½�v��ɣ��5���F�\�<;
�I�-GsK�#Y=s~H�D�'���q�����	��N˜k��]Q��r��yx��O�F��\���ǙK��?��$�W+�.�i�j�$���np}ś�t�aɏ�K#vĹE?�ۥvZN���~���
8�c����M_(n۱O��2oy̰�$�+h������h�)}:qĐA�*��/�	����3#�W+���@�Ԭ����
�A������8£q2�"��"�͏�?z4)x	�k�SO��]L? 3hH-�o�#�*�Y%���O�3��!@���,m[�SG��UN;I[��\Xѭ|�a�A�7�;x#Q�M,��b�s|�bYG�/O�*޲�������I�Ͳg=��|�kt$��ə�i礧"�gP�o&�ۯ���/R.��nG:��,���L�
fn�в�4Zs4
_�̲�\7yP��m��o��h|� ��A�W��@ �?Q|�%Ή��S�tH茺?�K(��9y�o���#�-��������:�Y@Vk���a���tM��[ɲ�
�T��{�ٹ��M��7F�\�4M`Lʂ{(&[IR;�PO��@:$�`�|_8K�M�ǳ��"PjQ� �C�l8��oܫ�$1�p�D�� ȵ����ˎ`�\p�1��-x3K8mǇ�"��覷��L���q�?�A�=��#�lTpOi[�K�Wn���v�V�K�ǔІ��X�b���!��l����Z=b��*BO�<jvS�`���YRt���]g%��;��@�w9Ro����.1���Â�d]*�+��6��� ���{�����RL����oW�Q�����Pd���UT�n�'�g�'p�4/s��Og[I'9~�rͻ�е�s�%��y��9r�ӏЭ8�C5Yu˵0і��J���4� h �C��+hoc�����`�����疴2�g*Lh,�?G� I�֖���~ܐ�8������0����0L)���;��W	�W��F3���I{	�N=�6*�^7`�d�Ɣ�盏������� ����q�k�J!�sm{B���Ǌ#��b
��	�Q8ʐ����lK����h��0	�+a�?hջ���9�M��>�8ߛ���1�<��-���gv!I�������4����æ������}��B��/\}�H��t��ؐ����k��L��˕t���e�t�6�S<)�8��У�U˰tc�5�Բ���堡yb���V9>n?�(��B��֧��`���N��}C=-�(��]j��G��0��&9H���P�4[�/�H�8�9�6�^���.i�Uɜ=������P�;݋ ����{H�^���j��Ĩ"�7�>}0�7��C��eTkk}ԝ����x/�;C�@c�TX�?kM[��T0ǘ�9l�ػ{��:%��joPI�� ߝ�D>�~�! �2� ^τU5� y��rA�) �.�I�k��gF� 2����ڠ"��Z5�a�3���6� ������ ;�X1��'_2�v���\_���yk�+#"{��8m'?2�;v1[k��~���a����Xt�w���׷44V��8�U7�z�9�£4G:k�X�m�/�Sω�D���}k�V�!�н�l���DF7�:�q�5̙�S�'As����z��f��J^#�!!9Wݦs:ꗜc[)eBf�:����v&Y'�%jU�,�bF�1��M%$�T���I����L�d6�l���-�8������0ؾ~b�juG�S�WMn9�^�dM�(�G�`'/��^&�,Sjӡ�T�b��,\���VX�(1�7|����ܖ�jx:�w���T[/a�5$�g�g{�l�\%�?˕p\]_�Z�����y c>@�T��I��eK���za~�@s>��"+)ESd��e������%H�L}�˄rV%+'��!=IM?��K[}B�+��p��ߍ�J��ݱi.����I��`�A#AJL:!�g�[�9����\� ��'����6^6�\`5j'�I�Mx�NDFD�n�M��Xe�7ހ�Z2/�@)D�����R�]�e��dp���*�F' �a045i?��2���h��P�l�`bP%
O�Oϕ�Y
�J�d��n�0���#Hfɤ�n4g��a�����|�*�|Shx�?��܈�z�t$ZK���AO(47�a����T|.C����@�����s���c�	��.���Č��;�x.�������pR��w�Osv�qCZ��{��o�A%�-6����+�t_)K8k���ʳs%YM�#ژw{S��b�:�AAa�mhWLĕ@�t\rTC��U/ԑ���1SsV?�M����fKAqh�ӝrFin�6xR��j�#9ʝz�ȍ1�Qk�� h�EJ�#B҅��J&��O�_'0/*���I�C���>�(�Q��To��	��1� �E����vo�]+��@��ˋ���'!"��-oG�Ø�[��7��ċ{��� 繽�|�<V�X~yk�p,��X T.�Gu���Y��W�����v��r����N��1�R��!y����il)|h�h�;�eؖy���v�ݨ];��\�Q_XY.ˊd-�R��g��gcݰ�K��9�V�.W��π�
u/"h�i3A��L���#�Xъ4��F~_`��(�)�P%�Ν�v���2��̾p��d�3���cql9(}J�B3�e�I�Y���t|]D=ӜcH�����#K ݃aP���A���,D�����Ɯj3����,1m'��M�p1�������y�K~�|[\U�������D�^,�_��PJ�-YZ�6b��IXv�B�d�]\Y��>�b���������nvߜ������v�s���#m�6z��Df�KĬ0VrO0_��Ź*�Ke�L$"�v*�1�a���H80~Ns8��1�O�?��E�LC�>�M�%&6��6�*���/u��c8I�z�Ur���8�<JG��i
�4�t7Ic�
�#_�-�z�ě�@��9�s>F�al�#�Ҝ�����jfnA��q��U=?��n�Q9z��Z.Z�E�q#�����:�xIa�<�wAM�����FBY��v�����;�OB�o{�ќ��R���XMO��E.8zo����yz������R}A�؂�$e�>_�F���9티�,4�~�N �a��oE�]�`�@��[Д�˅^@.	v�N�b��D��|Ы���"A\]�Z�E�E�-���r"U(QoW"���V�~�8�_,=b�����{G��[�l;4�~��-`���,�4�QRi����1��N?Qɣk�T,�M�<��J8v��D�Baih�tk"G�DU|���%]P�sX���@�uJ�h��4�_Ź;����D3�s��#�S������~Q^#1Y1NnX�x�u����PC����gi|\��WZ7绚�2-c ����JL���Ԙ����>�����<�������QJ	~�F˨���c�ހ�1�{��)�\)%�?���S�G͖��~f��W�:{�>��-��