��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�~�����tC�ޜ솚�*������Q鐙>��  �=C�B�~����/�kt��*��x�KN����Dʱ9]
����tW��2S;c�jZc{�?��!b�$^��[v��W,�ީ��+O�N\L��B�!t�XE�"C �n��˾�w�,C6�nSb�N��t� t�';��\/�X`��.�ó[�g��8!�� ߪZ敁��ļ��ۺ$3���m]Z��7;!�՟£��z��u�.��W����9�	����	�a�Q���߆��)�O3{��f��$���!�rq۬��"�<��"Ӄ���b�0U����I��W�_An��Mz�d_���K��w�7�MnPe{*����������.Xb
�=��9݃i���|�'�$U���{�Q�z�.c���:��1j��S���{��*_�zwȀC�D���J�"�
�F��C�����mq�]��d����Q�pYgك����&��f_� �!IكZ���=��|Z�f��b��,=xV0O#y�[|� 1jB�sg�Z�݇�5�~��;��U=��w�aB��ao��4k�[���*���v��GF�xe�v������^�1��R!O�!L��<N����tj��� �)Z2��}��$�>�Gk�p��-�,�Lm��n���Jۉ5V􂘉�d#���!��XQQ}s��Hw��j�e��7�B�Rt�t���VInd�Q،w�/���I��晼��>����_�/x������f�ƿ�uH��hߝm�)��4���N�:d�^k��e���N��4��F������l.��� Ps淼���s�����:/@�X^ԭ%���'-�x�G*�vY���3�W�/�%�����xq �N���:n�'4_�B����b��$l�u��|�w��lH�sh��+Dv
���u����u����������s�ѓ����w�õ6
~[[�C��u�f|����/&\4rCR!� UZ[�ۻu쎽��[o�v�Ho[g*$�`�dX������b��wT��%?��\q��^TP�š�5n/>%����a�8_!����'wC�p�)��a!�����h���Q��7�ȡ�g\�]rގj���ޔqb�HV�z	/�!��ev�*��I.��!�P��&XD���)�bY�7�X�aC.��=ac��P�>(�P�.�H�~[0!���O��򹷌5D���	;! Ͷ`�(��M�FY�g�5�!(L�:��)�S����9$o�3"Sub�/�u�1��%�L!��T?�$��[��w.���.�CX�A_����-.��D�l^l\�z{,��7�{�J��Ӭ����yb~j-�tp�`����� ��G���2��_�g��6Lj�>!���V@�k"�U���PwD�L�Q��pϞj	h�d�6Zs8Y�D{{�s*}���/�O����.[j(K�)�)�#0pZ��Qd�2=�X6����b2��wo��Z�E��3�k���d�(ڝ�_�D&l��)��e���L��6E���^���x���kfԟ|m�A�P�0a�;�A���]��"Ă!�x#{W�4,��dǿ1 Y"�:27qu8Gܧ��9v�+��J�4��G~�"�4?�up�qe�9s%���R����R��PZ4���!���)��艹hh�D��KW7rp8ύW2�5u��>�k1 ��Bd���wX��/�����zͲ����m�o=��A����-� �R� ��Ԇ%o��`_a��}C̫��o���t>.3� ���EP�a��4�U�í�� Y�Q���cz	0|����Ne�������z��Zt��4U���tl��t��f�`Lw�Z�i7�wN��M?�@�Jk��?�
3�3l!��*�*��Cex���hwj^%ۅݛ�4���R��H�j���Ķ�}og=NV�&i3���2S��	��`z��V��	qP�����)f�Z�V����_��O"�}����]���iG�)�<����ې��+��eo/(JvO����t�ؘ���s=K��t_ھ�k�3U����r�����#��1뻋�m���گ�v���|�䗜!�|m�*w?��m�7ĺH˾���E�����4�r��8��-�ʃ"�����e�{�+=�:�2��0�������Q��S�p-�v/�BK�*ݷ��_�i~ē�0u3���&��{ݰ��U����O⠨펼��}]�/��vk�X<ܠ�X=iY��rhh�v%��i���� $�B[ZNJ'D���x0'�z��m�%����oT~�㪨�	/�(����1�HYH��X���_�#a�tu2�.���6|��9b�`��6�_o�lvk�""bK00��'��aC��)�|�GТ��v��2�,�r���V�9ޢkK���.,*�+����Z�Ҧ�7E�s% �y�*t�p��֡�saӳ�jE�]Q���=�[e?�$��,;lVU�8lk�`��j,r���t���y�s��e�J�ó�Z[�-���Fj�g`z׼"�X��O�Դ�����g�"�����s�\F��ᮊ��J��S��H�dJ;h3J�ԓ:�"�>��.6 N�>@�3c�߸�Co�'C����>�FL��vuUҞN41.�X���=幥�Tזg�hAW�4�l�2��ɽ<�)����*V�J� ��;2�V �	����D�?YҌ��1��@am�vw%�P%cG�;9�k�P��R,58m�U���n���@~:�v�qS(�f�v��b��w�Q����m j��]G�?#�X�C�>�1?�6_�Ҧu��Ġ��@;����=���¾|�Z������ ���V����>���:��;�֍��AM����9����X�����oS��G.��"L�����_���(�e�A��2&�CJ��5�Mn�f'x��͐>�V�]����J��F��4���@�n�VT�����%q������x�	m���jUIO݋���H�6����[����V�U���3�P�7�g��sd���'���j�<F��q�m��,s��=�F�k#@~��s7G�/xҭ+�Z�(%�x�WR��|�(Ԑ'-OR�PnZ�ry`a.,�w2�}�X�e+�d�]%��*����DLgq�ȁ6]%.�v�B��
�^z�}T̩�cu��;��q�	�NY�U�\ޭ����`"=eI=�&�s��t+��2e����q�w�C�>�#�Z�Z��Dg�>�"TSAڑ��A��v��]�0r�2�����:�����kx�B�R��s|�eֵ]�{Q��=���g�|�#(�ܐ�O*	�8��g�.��o�O�������Zn���/#՟��h����v]���x����%�o�'z��1�v�j�$)>R�[w��S�w��qƳ�.�q�9�-���-X��4sf���'�D&�[�*�5��ˇ���;���ݩ%����Ec�Ҕ��tTip2��Vw�sS󝾍QAz�ة&�q��Tpt�L��>V������c|RW��21�Ҧ�`�I�@�(`�8֗oG���|#�T�����pf�`�����GP`Z��&���ȊY����8r}�}�s��!V�C�J�]���K)���P.$�}A5-��Z������8�P�#��x��:}T�l��mC?�:��݋Gܪ����#��(���>�D�:���dQ0YQ�2�E�9EP[,���xӞv����tب���-�d1�x@�<�fMè��	�)-�	�NL�����d�AC9��4ya5
of��M�Z�Z~c�k!�+:��k���m(�6?�y��u���P�����I�G?��U�D�1PE�{!Z2#�k���j~��omKؑ�R�N�ɣ��j����	~>����=_��b�v��L^K(�Ե���������59�?E�#��X��O~'����>��,��i'i���܌�bk�<;C:�l9W����T"i^��ڮ�V���+(�zp=��<Y*�N<��k��!���;�,߇���b�|�'h��ڞ����ω�6�Ԙ�t%�:J8�j���fx:u�q��2�T\����^���%�R��X�N��B����X%}8���Y�ܢ7�L