��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�_#jo��a�>�)B����IB�m
��.�E3^������rLx�"�`g�!9O#�����,��眽J�����"�Q�|7�e��v(<J�h�&�" ��y;$�G�6ը���'�}�K���nN�H!��W��@� �c�f��i~��|"ޟ�Ѱ���;�W#h�0%�37}EOΤ�#��B������l}��mG���M2�:�Ld�B�k(�T��LG����5>zA/I��T��Z���1%|D)F��R���r���5�'�i��+�Xz3W��|��_ŵ|�%(�T-$��(�>�L^y�_�W�/�V�4���,Wn,��ɻ��WO�p��H����� �	��'gm[�� C'"\&\F�82�C{c�&6h-�0.�N�����M#i�6b�[�@�ʹY����|��-O�����P^�]~ju�c�=`�[���$ɍ�k�r~ֻf&U�[��\F	*��gG�5���vC"�ۨX���z��c�����
K����D=�����qv�8D)������;�,/�ȃ�
�A�kM���[�,�ikY/l	o��G�/��8&RdFt"��y������0c����|�X&ç�E�>%�z���kz�@]�$��O��O��F�y>F�%h�x��~��5.