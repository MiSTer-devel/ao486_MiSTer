// system.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_clk,             //        clk.clk
		output wire        clk_sys_clk,         //    clk_sys.clk
		input  wire        cpu_reset_reset,     //  cpu_reset.reset
		output wire [31:0] ddram_address,       //      ddram.address
		output wire        ddram_read,          //           .read
		input  wire        ddram_waitrequest,   //           .waitrequest
		input  wire [63:0] ddram_readdata,      //           .readdata
		output wire        ddram_write,         //           .write
		output wire [63:0] ddram_writedata,     //           .writedata
		input  wire        ddram_readdatavalid, //           .readdatavalid
		output wire [7:0]  ddram_byteenable,    //           .byteenable
		output wire [7:0]  ddram_burstcount,    //           .burstcount
		output wire        disk_op_read,        //       disk.op_read
		output wire        disk_op_write,       //           .op_write
		input  wire        disk_result_ok,      //           .result_ok
		input  wire        disk_result_error,   //           .result_error
		output wire        disk_op_device,      //           .op_device
		output wire        mem_waitrequest,     //        mem.waitrequest
		output wire [31:0] mem_readdata,        //           .readdata
		output wire        mem_readdatavalid,   //           .readdatavalid
		input  wire [0:0]  mem_burstcount,      //           .burstcount
		input  wire [31:0] mem_writedata,       //           .writedata
		input  wire [31:0] mem_address,         //           .address
		input  wire        mem_write,           //           .write
		input  wire        mem_read,            //           .read
		input  wire [3:0]  mem_byteenable,      //           .byteenable
		input  wire        mem_debugaccess,     //           .debugaccess
		input  wire        pll_reset_reset,     //  pll_reset.reset
		input  wire        ps2_kbclk_in,        //        ps2.kbclk_in
		input  wire        ps2_kbdat_in,        //           .kbdat_in
		output wire        ps2_kbclk_out,       //           .kbclk_out
		output wire        ps2_kbdat_out,       //           .kbdat_out
		input  wire        ps2_mouseclk_in,     //           .mouseclk_in
		input  wire        ps2_mousedat_in,     //           .mousedat_in
		output wire        ps2_mouseclk_out,    //           .mouseclk_out
		output wire        ps2_mousedat_out,    //           .mousedat_out
		output wire        ps2_misc_a20_enable, //   ps2_misc.a20_enable
		output wire        ps2_misc_reset_n,    //           .reset_n
		input  wire        qsys_reset_reset,    // qsys_reset.reset
		output wire [15:0] sound_sample_l,      //      sound.sample_l
		output wire [15:0] sound_sample_r,      //           .sample_r
		input  wire        sound_fm_mode,       //           .fm_mode
		input  wire        sound_mpu_midi_in,   //           .mpu_midi_in
		output wire        sound_mpu_midi_out,  //           .mpu_midi_out
		output wire        speaker_enable,      //    speaker.enable
		output wire        speaker_out,         //           .out
		input  wire        uart_h_cts_n,        //     uart_h.cts_n
		output wire        uart_h_rts_n,        //           .rts_n
		input  wire        uart_h_dsr_n,        //           .dsr_n
		input  wire        uart_h_dcd_n,        //           .dcd_n
		input  wire        uart_h_ri_n,         //           .ri_n
		output wire        uart_h_dtr_n,        //           .dtr_n
		output wire        uart_h_out1_n,       //           .out1_n
		output wire        uart_h_out2_n,       //           .out2_n
		input  wire        uart_s_sin,          //     uart_s.sin
		output wire        uart_s_sout,         //           .sout
		output wire        uart_s_sout_oe,      //           .sout_oe
		output wire        vga_clock,           //        vga.clock
		output wire        vga_blank_n,         //           .blank_n
		output wire        vga_hsync,           //           .hsync
		output wire        vga_vsync,           //           .vsync
		output wire [7:0]  vga_r,               //           .r
		output wire [7:0]  vga_g,               //           .g
		output wire [7:0]  vga_b                //           .b
	);

	wire         ao486_avalon_memory_waitrequest;                                      // pc_bus:mem_waitrequest -> ao486:avm_waitrequest
	wire  [31:0] ao486_avalon_memory_readdata;                                         // pc_bus:mem_readdata -> ao486:avm_readdata
	wire  [29:0] ao486_avalon_memory_address;                                          // ao486:avm_address -> pc_bus:mem_address
	wire   [3:0] ao486_avalon_memory_byteenable;                                       // ao486:avm_byteenable -> pc_bus:mem_byteenable
	wire         ao486_avalon_memory_read;                                             // ao486:avm_read -> pc_bus:mem_read
	wire         ao486_avalon_memory_readdatavalid;                                    // pc_bus:mem_readdatavalid -> ao486:avm_readdatavalid
	wire  [31:0] ao486_avalon_memory_writedata;                                        // ao486:avm_writedata -> pc_bus:mem_writedata
	wire         ao486_avalon_memory_write;                                            // ao486:avm_write -> pc_bus:mem_write
	wire   [2:0] ao486_avalon_memory_burstcount;                                       // ao486:avm_burstcount -> pc_bus:mem_burstcount
	wire  [31:0] width_trans_out_readdata;                                             // uart:readdata -> width_trans:out_readdata
	wire   [8:0] width_trans_out_address;                                              // width_trans:out_address -> uart:addr
	wire         width_trans_out_read;                                                 // width_trans:out_read -> uart:read
	wire         width_trans_out_write;                                                // width_trans:out_write -> uart:write
	wire  [31:0] width_trans_out_writedata;                                            // width_trans:out_writedata -> uart:writedata
	wire         pll_0_outclk1_clk;                                                    // pll_0:outclk_1 -> vga:clk_vga
	wire         pll_0_outclk2_clk;                                                    // pll_0:outclk_2 -> [irq_synchronizer:receiver_clk, mm_interconnect_0:pll_0_outclk2_clk, rst_controller_001:clk, uart:clk, width_trans:clk]
	wire         ps2_conduit_a20_a20_enable;                                           // ps2:a20_enable -> ao486:a20_enable
	wire   [7:0] pc_dma_conduit_dma_floppy_dma_floppy_readdata;                        // pc_dma:dma_floppy_readdata -> floppy0:dma_floppy_readdata
	wire         pc_dma_conduit_dma_floppy_dma_floppy_terminal;                        // pc_dma:dma_floppy_terminal -> floppy0:dma_floppy_terminal
	wire   [7:0] floppy0_conduit_dma_floppy_dma_floppy_writedata;                      // floppy0:dma_floppy_writedata -> pc_dma:dma_floppy_writedata
	wire         floppy0_conduit_dma_floppy_dma_floppy_req;                            // floppy0:dma_floppy_req -> pc_dma:dma_floppy_req
	wire         pc_dma_conduit_dma_floppy_dma_floppy_ack;                             // pc_dma:dma_floppy_ack -> floppy0:dma_floppy_ack
	wire         sound_conduit_dma_soundblaster_dma_soundblaster_req;                  // sound:dma_soundblaster_req -> pc_dma:dma_soundblaster_req
	wire         pc_dma_conduit_dma_soundblaster_dma_soundblaster_terminal;            // pc_dma:dma_soundblaster_terminal -> sound:dma_soundblaster_terminal
	wire   [7:0] pc_dma_conduit_dma_soundblaster_dma_soundblaster_readdata;            // pc_dma:dma_soundblaster_readdata -> sound:dma_soundblaster_readdata
	wire   [7:0] sound_conduit_dma_soundblaster_dma_soundblaster_writedata;            // sound:dma_soundblaster_writedata -> pc_dma:dma_soundblaster_writedata
	wire         pc_dma_conduit_dma_soundblaster_dma_soundblaster_ack;                 // pc_dma:dma_soundblaster_ack -> sound:dma_soundblaster_ack
	wire   [7:0] hdd0_conduit_ide_3f6_ide_3f6_readdata;                                // hdd0:ide_3f6_readdata -> floppy0:ide_3f6_readdata
	wire   [7:0] floppy0_conduit_ide_3f6_ide_3f6_writedata;                            // floppy0:ide_3f6_writedata -> hdd0:ide_3f6_writedata
	wire         floppy0_conduit_ide_3f6_ide_3f6_write;                                // floppy0:ide_3f6_write -> hdd0:ide_3f6_write
	wire         floppy0_conduit_ide_3f6_ide_3f6_read;                                 // floppy0:ide_3f6_read -> hdd0:ide_3f6_read
	wire   [7:0] hdd1_conduit_ide_3f6_ide_3f6_readdata;                                // hdd1:ide_3f6_readdata -> hddext_0x370:ide_3f6_readdata
	wire   [7:0] hddext_0x370_conduit_ide_3f6_ide_3f6_writedata;                       // hddext_0x370:ide_3f6_writedata -> hdd1:ide_3f6_writedata
	wire         hddext_0x370_conduit_ide_3f6_ide_3f6_write;                           // hddext_0x370:ide_3f6_write -> hdd1:ide_3f6_write
	wire         hddext_0x370_conduit_ide_3f6_ide_3f6_read;                            // hddext_0x370:ide_3f6_read -> hdd1:ide_3f6_read
	wire         ao486_interrupt_interrupt_done;                                       // ao486:interrupt_done -> pic:interrupt_done
	wire         pic_conduit_interrupt_interrupt_do;                                   // pic:interrupt_do -> ao486:interrupt_do
	wire   [7:0] pic_conduit_interrupt_interrupt_vector;                               // pic:interrupt_vector -> ao486:interrupt_vector
	wire         ps2_conduit_speaker_61h_speaker_61h_read;                             // ps2:speaker_61h_read -> pit:speaker_61h_read
	wire         ps2_conduit_speaker_61h_speaker_61h_write;                            // ps2:speaker_61h_write -> pit:speaker_61h_write
	wire   [7:0] pit_conduit_speaker_61h_speaker_61h_readdata;                         // pit:speaker_61h_readdata -> ps2:speaker_61h_readdata
	wire   [7:0] ps2_conduit_speaker_61h_speaker_61h_writedata;                        // ps2:speaker_61h_writedata -> pit:speaker_61h_writedata
	wire         reset_sys_reset_out_reset;                                            // reset_sys:reset_out -> [address_span_extender:reset, driver_sd:rst_n, floppy0:rst_n, hdd0:rst_n, hdd1:rst_n, hddext_0x370:rst_n, irq_mapper:reset, irq_synchronizer:sender_reset, mm_bridge:reset, mm_interconnect_0:sound_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:floppy0_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_3:pc_bus_reset_sink_reset_bridge_in_reset_reset, pc_bus:rst_n, pc_dma:rst_n, pic:rst_n, pit:rst_n, ps2:rst_n, rst_controller_001:reset_in0, rtc:rst_n, sound:rst_n, vga:rst_n]
	wire  [31:0] ao486_avalon_io_readdata;                                             // mm_interconnect_0:ao486_avalon_io_readdata -> ao486:avalon_io_readdata
	wire         ao486_avalon_io_waitrequest;                                          // mm_interconnect_0:ao486_avalon_io_waitrequest -> ao486:avalon_io_waitrequest
	wire  [15:0] ao486_avalon_io_address;                                              // ao486:avalon_io_address -> mm_interconnect_0:ao486_avalon_io_address
	wire   [3:0] ao486_avalon_io_byteenable;                                           // ao486:avalon_io_byteenable -> mm_interconnect_0:ao486_avalon_io_byteenable
	wire         ao486_avalon_io_read;                                                 // ao486:avalon_io_read -> mm_interconnect_0:ao486_avalon_io_read
	wire         ao486_avalon_io_readdatavalid;                                        // mm_interconnect_0:ao486_avalon_io_readdatavalid -> ao486:avalon_io_readdatavalid
	wire         ao486_avalon_io_write;                                                // ao486:avalon_io_write -> mm_interconnect_0:ao486_avalon_io_write
	wire  [31:0] ao486_avalon_io_writedata;                                            // ao486:avalon_io_writedata -> mm_interconnect_0:ao486_avalon_io_writedata
	wire   [7:0] mm_interconnect_0_sound_fm_readdata;                                  // sound:fm_readdata -> mm_interconnect_0:sound_fm_readdata
	wire   [1:0] mm_interconnect_0_sound_fm_address;                                   // mm_interconnect_0:sound_fm_address -> sound:fm_address
	wire         mm_interconnect_0_sound_fm_read;                                      // mm_interconnect_0:sound_fm_read -> sound:fm_read
	wire         mm_interconnect_0_sound_fm_write;                                     // mm_interconnect_0:sound_fm_write -> sound:fm_write
	wire   [7:0] mm_interconnect_0_sound_fm_writedata;                                 // mm_interconnect_0:sound_fm_writedata -> sound:fm_writedata
	wire   [7:0] mm_interconnect_0_width_trans_in_readdata;                            // width_trans:in_readdata -> mm_interconnect_0:width_trans_in_readdata
	wire   [2:0] mm_interconnect_0_width_trans_in_address;                             // mm_interconnect_0:width_trans_in_address -> width_trans:in_address
	wire         mm_interconnect_0_width_trans_in_read;                                // mm_interconnect_0:width_trans_in_read -> width_trans:in_read
	wire         mm_interconnect_0_width_trans_in_write;                               // mm_interconnect_0:width_trans_in_write -> width_trans:in_write
	wire   [7:0] mm_interconnect_0_width_trans_in_writedata;                           // mm_interconnect_0:width_trans_in_writedata -> width_trans:in_writedata
	wire   [7:0] mm_interconnect_0_sound_io_readdata;                                  // sound:io_readdata -> mm_interconnect_0:sound_io_readdata
	wire   [3:0] mm_interconnect_0_sound_io_address;                                   // mm_interconnect_0:sound_io_address -> sound:io_address
	wire         mm_interconnect_0_sound_io_read;                                      // mm_interconnect_0:sound_io_read -> sound:io_read
	wire         mm_interconnect_0_sound_io_write;                                     // mm_interconnect_0:sound_io_write -> sound:io_write
	wire   [7:0] mm_interconnect_0_sound_io_writedata;                                 // mm_interconnect_0:sound_io_writedata -> sound:io_writedata
	wire   [7:0] mm_interconnect_0_rtc_io_readdata;                                    // rtc:io_readdata -> mm_interconnect_0:rtc_io_readdata
	wire   [0:0] mm_interconnect_0_rtc_io_address;                                     // mm_interconnect_0:rtc_io_address -> rtc:io_address
	wire         mm_interconnect_0_rtc_io_read;                                        // mm_interconnect_0:rtc_io_read -> rtc:io_read
	wire         mm_interconnect_0_rtc_io_write;                                       // mm_interconnect_0:rtc_io_write -> rtc:io_write
	wire   [7:0] mm_interconnect_0_rtc_io_writedata;                                   // mm_interconnect_0:rtc_io_writedata -> rtc:io_writedata
	wire   [7:0] mm_interconnect_0_pit_io_readdata;                                    // pit:io_readdata -> mm_interconnect_0:pit_io_readdata
	wire   [1:0] mm_interconnect_0_pit_io_address;                                     // mm_interconnect_0:pit_io_address -> pit:io_address
	wire         mm_interconnect_0_pit_io_read;                                        // mm_interconnect_0:pit_io_read -> pit:io_read
	wire         mm_interconnect_0_pit_io_write;                                       // mm_interconnect_0:pit_io_write -> pit:io_write
	wire   [7:0] mm_interconnect_0_pit_io_writedata;                                   // mm_interconnect_0:pit_io_writedata -> pit:io_writedata
	wire  [31:0] mm_interconnect_0_hdd0_io_readdata;                                   // hdd0:io_readdata -> mm_interconnect_0:hdd0_io_readdata
	wire   [0:0] mm_interconnect_0_hdd0_io_address;                                    // mm_interconnect_0:hdd0_io_address -> hdd0:io_address
	wire         mm_interconnect_0_hdd0_io_read;                                       // mm_interconnect_0:hdd0_io_read -> hdd0:io_read
	wire   [3:0] mm_interconnect_0_hdd0_io_byteenable;                                 // mm_interconnect_0:hdd0_io_byteenable -> hdd0:io_byteenable
	wire         mm_interconnect_0_hdd0_io_write;                                      // mm_interconnect_0:hdd0_io_write -> hdd0:io_write
	wire  [31:0] mm_interconnect_0_hdd0_io_writedata;                                  // mm_interconnect_0:hdd0_io_writedata -> hdd0:io_writedata
	wire   [7:0] mm_interconnect_0_floppy0_io_readdata;                                // floppy0:io_readdata -> mm_interconnect_0:floppy0_io_readdata
	wire   [2:0] mm_interconnect_0_floppy0_io_address;                                 // mm_interconnect_0:floppy0_io_address -> floppy0:io_address
	wire         mm_interconnect_0_floppy0_io_read;                                    // mm_interconnect_0:floppy0_io_read -> floppy0:io_read
	wire         mm_interconnect_0_floppy0_io_write;                                   // mm_interconnect_0:floppy0_io_write -> floppy0:io_write
	wire   [7:0] mm_interconnect_0_floppy0_io_writedata;                               // mm_interconnect_0:floppy0_io_writedata -> floppy0:io_writedata
	wire   [7:0] mm_interconnect_0_ps2_io_readdata;                                    // ps2:io_readdata -> mm_interconnect_0:ps2_io_readdata
	wire   [2:0] mm_interconnect_0_ps2_io_address;                                     // mm_interconnect_0:ps2_io_address -> ps2:io_address
	wire         mm_interconnect_0_ps2_io_read;                                        // mm_interconnect_0:ps2_io_read -> ps2:io_read
	wire         mm_interconnect_0_ps2_io_write;                                       // mm_interconnect_0:ps2_io_write -> ps2:io_write
	wire   [7:0] mm_interconnect_0_ps2_io_writedata;                                   // mm_interconnect_0:ps2_io_writedata -> ps2:io_writedata
	wire  [31:0] mm_interconnect_0_hdd1_io_readdata;                                   // hdd1:io_readdata -> mm_interconnect_0:hdd1_io_readdata
	wire   [0:0] mm_interconnect_0_hdd1_io_address;                                    // mm_interconnect_0:hdd1_io_address -> hdd1:io_address
	wire         mm_interconnect_0_hdd1_io_read;                                       // mm_interconnect_0:hdd1_io_read -> hdd1:io_read
	wire   [3:0] mm_interconnect_0_hdd1_io_byteenable;                                 // mm_interconnect_0:hdd1_io_byteenable -> hdd1:io_byteenable
	wire         mm_interconnect_0_hdd1_io_write;                                      // mm_interconnect_0:hdd1_io_write -> hdd1:io_write
	wire  [31:0] mm_interconnect_0_hdd1_io_writedata;                                  // mm_interconnect_0:hdd1_io_writedata -> hdd1:io_writedata
	wire   [7:0] mm_interconnect_0_hddext_0x370_io_readdata;                           // hddext_0x370:io_readdata -> mm_interconnect_0:hddext_0x370_io_readdata
	wire   [2:0] mm_interconnect_0_hddext_0x370_io_address;                            // mm_interconnect_0:hddext_0x370_io_address -> hddext_0x370:io_address
	wire         mm_interconnect_0_hddext_0x370_io_read;                               // mm_interconnect_0:hddext_0x370_io_read -> hddext_0x370:io_read
	wire         mm_interconnect_0_hddext_0x370_io_write;                              // mm_interconnect_0:hddext_0x370_io_write -> hddext_0x370:io_write
	wire   [7:0] mm_interconnect_0_hddext_0x370_io_writedata;                          // mm_interconnect_0:hddext_0x370_io_writedata -> hddext_0x370:io_writedata
	wire   [7:0] mm_interconnect_0_vga_io_b_readdata;                                  // vga:io_b_readdata -> mm_interconnect_0:vga_io_b_readdata
	wire   [3:0] mm_interconnect_0_vga_io_b_address;                                   // mm_interconnect_0:vga_io_b_address -> vga:io_b_address
	wire         mm_interconnect_0_vga_io_b_read;                                      // mm_interconnect_0:vga_io_b_read -> vga:io_b_read
	wire         mm_interconnect_0_vga_io_b_write;                                     // mm_interconnect_0:vga_io_b_write -> vga:io_b_write
	wire   [7:0] mm_interconnect_0_vga_io_b_writedata;                                 // mm_interconnect_0:vga_io_b_writedata -> vga:io_b_writedata
	wire   [7:0] mm_interconnect_0_vga_io_c_readdata;                                  // vga:io_c_readdata -> mm_interconnect_0:vga_io_c_readdata
	wire   [3:0] mm_interconnect_0_vga_io_c_address;                                   // mm_interconnect_0:vga_io_c_address -> vga:io_c_address
	wire         mm_interconnect_0_vga_io_c_read;                                      // mm_interconnect_0:vga_io_c_read -> vga:io_c_read
	wire         mm_interconnect_0_vga_io_c_write;                                     // mm_interconnect_0:vga_io_c_write -> vga:io_c_write
	wire   [7:0] mm_interconnect_0_vga_io_c_writedata;                                 // mm_interconnect_0:vga_io_c_writedata -> vga:io_c_writedata
	wire   [7:0] mm_interconnect_0_vga_io_d_readdata;                                  // vga:io_d_readdata -> mm_interconnect_0:vga_io_d_readdata
	wire   [3:0] mm_interconnect_0_vga_io_d_address;                                   // mm_interconnect_0:vga_io_d_address -> vga:io_d_address
	wire         mm_interconnect_0_vga_io_d_read;                                      // mm_interconnect_0:vga_io_d_read -> vga:io_d_read
	wire         mm_interconnect_0_vga_io_d_write;                                     // mm_interconnect_0:vga_io_d_write -> vga:io_d_write
	wire   [7:0] mm_interconnect_0_vga_io_d_writedata;                                 // mm_interconnect_0:vga_io_d_writedata -> vga:io_d_writedata
	wire   [7:0] mm_interconnect_0_pc_dma_master_readdata;                             // pc_dma:master_readdata -> mm_interconnect_0:pc_dma_master_readdata
	wire   [4:0] mm_interconnect_0_pc_dma_master_address;                              // mm_interconnect_0:pc_dma_master_address -> pc_dma:master_address
	wire         mm_interconnect_0_pc_dma_master_read;                                 // mm_interconnect_0:pc_dma_master_read -> pc_dma:master_read
	wire         mm_interconnect_0_pc_dma_master_write;                                // mm_interconnect_0:pc_dma_master_write -> pc_dma:master_write
	wire   [7:0] mm_interconnect_0_pc_dma_master_writedata;                            // mm_interconnect_0:pc_dma_master_writedata -> pc_dma:master_writedata
	wire   [7:0] mm_interconnect_0_pic_master_readdata;                                // pic:master_readdata -> mm_interconnect_0:pic_master_readdata
	wire   [0:0] mm_interconnect_0_pic_master_address;                                 // mm_interconnect_0:pic_master_address -> pic:master_address
	wire         mm_interconnect_0_pic_master_read;                                    // mm_interconnect_0:pic_master_read -> pic:master_read
	wire         mm_interconnect_0_pic_master_write;                                   // mm_interconnect_0:pic_master_write -> pic:master_write
	wire   [7:0] mm_interconnect_0_pic_master_writedata;                               // mm_interconnect_0:pic_master_writedata -> pic:master_writedata
	wire   [7:0] mm_interconnect_0_sound_mpu_readdata;                                 // sound:mpu_readdata -> mm_interconnect_0:sound_mpu_readdata
	wire   [2:0] mm_interconnect_0_sound_mpu_address;                                  // mm_interconnect_0:sound_mpu_address -> sound:mpu_address
	wire         mm_interconnect_0_sound_mpu_read;                                     // mm_interconnect_0:sound_mpu_read -> sound:mpu_read
	wire         mm_interconnect_0_sound_mpu_write;                                    // mm_interconnect_0:sound_mpu_write -> sound:mpu_write
	wire   [7:0] mm_interconnect_0_sound_mpu_writedata;                                // mm_interconnect_0:sound_mpu_writedata -> sound:mpu_writedata
	wire   [7:0] mm_interconnect_0_pc_dma_page_readdata;                               // pc_dma:page_readdata -> mm_interconnect_0:pc_dma_page_readdata
	wire   [3:0] mm_interconnect_0_pc_dma_page_address;                                // mm_interconnect_0:pc_dma_page_address -> pc_dma:page_address
	wire         mm_interconnect_0_pc_dma_page_read;                                   // mm_interconnect_0:pc_dma_page_read -> pc_dma:page_read
	wire         mm_interconnect_0_pc_dma_page_write;                                  // mm_interconnect_0:pc_dma_page_write -> pc_dma:page_write
	wire   [7:0] mm_interconnect_0_pc_dma_page_writedata;                              // mm_interconnect_0:pc_dma_page_writedata -> pc_dma:page_writedata
	wire   [7:0] mm_interconnect_0_pc_dma_slave_readdata;                              // pc_dma:slave_readdata -> mm_interconnect_0:pc_dma_slave_readdata
	wire   [3:0] mm_interconnect_0_pc_dma_slave_address;                               // mm_interconnect_0:pc_dma_slave_address -> pc_dma:slave_address
	wire         mm_interconnect_0_pc_dma_slave_read;                                  // mm_interconnect_0:pc_dma_slave_read -> pc_dma:slave_read
	wire         mm_interconnect_0_pc_dma_slave_write;                                 // mm_interconnect_0:pc_dma_slave_write -> pc_dma:slave_write
	wire   [7:0] mm_interconnect_0_pc_dma_slave_writedata;                             // mm_interconnect_0:pc_dma_slave_writedata -> pc_dma:slave_writedata
	wire   [7:0] mm_interconnect_0_pic_slave_readdata;                                 // pic:slave_readdata -> mm_interconnect_0:pic_slave_readdata
	wire   [0:0] mm_interconnect_0_pic_slave_address;                                  // mm_interconnect_0:pic_slave_address -> pic:slave_address
	wire         mm_interconnect_0_pic_slave_read;                                     // mm_interconnect_0:pic_slave_read -> pic:slave_read
	wire         mm_interconnect_0_pic_slave_write;                                    // mm_interconnect_0:pic_slave_write -> pic:slave_write
	wire   [7:0] mm_interconnect_0_pic_slave_writedata;                                // mm_interconnect_0:pic_slave_writedata -> pic:slave_writedata
	wire   [7:0] mm_interconnect_0_ps2_sysctl_readdata;                                // ps2:sysctl_readdata -> mm_interconnect_0:ps2_sysctl_readdata
	wire   [3:0] mm_interconnect_0_ps2_sysctl_address;                                 // mm_interconnect_0:ps2_sysctl_address -> ps2:sysctl_address
	wire         mm_interconnect_0_ps2_sysctl_read;                                    // mm_interconnect_0:ps2_sysctl_read -> ps2:sysctl_read
	wire         mm_interconnect_0_ps2_sysctl_write;                                   // mm_interconnect_0:ps2_sysctl_write -> ps2:sysctl_write
	wire   [7:0] mm_interconnect_0_ps2_sysctl_writedata;                               // mm_interconnect_0:ps2_sysctl_writedata -> ps2:sysctl_writedata
	wire         floppy0_avalon_master_waitrequest;                                    // mm_interconnect_1:floppy0_avalon_master_waitrequest -> floppy0:sd_master_waitrequest
	wire  [31:0] floppy0_avalon_master_readdata;                                       // mm_interconnect_1:floppy0_avalon_master_readdata -> floppy0:sd_master_readdata
	wire  [31:0] floppy0_avalon_master_address;                                        // floppy0:sd_master_address -> mm_interconnect_1:floppy0_avalon_master_address
	wire         floppy0_avalon_master_read;                                           // floppy0:sd_master_read -> mm_interconnect_1:floppy0_avalon_master_read
	wire         floppy0_avalon_master_readdatavalid;                                  // mm_interconnect_1:floppy0_avalon_master_readdatavalid -> floppy0:sd_master_readdatavalid
	wire         floppy0_avalon_master_write;                                          // floppy0:sd_master_write -> mm_interconnect_1:floppy0_avalon_master_write
	wire  [31:0] floppy0_avalon_master_writedata;                                      // floppy0:sd_master_writedata -> mm_interconnect_1:floppy0_avalon_master_writedata
	wire         hdd0_avalon_master_waitrequest;                                       // mm_interconnect_1:hdd0_avalon_master_waitrequest -> hdd0:sd_master_waitrequest
	wire  [31:0] hdd0_avalon_master_readdata;                                          // mm_interconnect_1:hdd0_avalon_master_readdata -> hdd0:sd_master_readdata
	wire  [31:0] hdd0_avalon_master_address;                                           // hdd0:sd_master_address -> mm_interconnect_1:hdd0_avalon_master_address
	wire         hdd0_avalon_master_read;                                              // hdd0:sd_master_read -> mm_interconnect_1:hdd0_avalon_master_read
	wire         hdd0_avalon_master_readdatavalid;                                     // mm_interconnect_1:hdd0_avalon_master_readdatavalid -> hdd0:sd_master_readdatavalid
	wire         hdd0_avalon_master_write;                                             // hdd0:sd_master_write -> mm_interconnect_1:hdd0_avalon_master_write
	wire  [31:0] hdd0_avalon_master_writedata;                                         // hdd0:sd_master_writedata -> mm_interconnect_1:hdd0_avalon_master_writedata
	wire         hdd1_avalon_master_waitrequest;                                       // mm_interconnect_1:hdd1_avalon_master_waitrequest -> hdd1:sd_master_waitrequest
	wire  [31:0] hdd1_avalon_master_readdata;                                          // mm_interconnect_1:hdd1_avalon_master_readdata -> hdd1:sd_master_readdata
	wire  [31:0] hdd1_avalon_master_address;                                           // hdd1:sd_master_address -> mm_interconnect_1:hdd1_avalon_master_address
	wire         hdd1_avalon_master_read;                                              // hdd1:sd_master_read -> mm_interconnect_1:hdd1_avalon_master_read
	wire         hdd1_avalon_master_readdatavalid;                                     // mm_interconnect_1:hdd1_avalon_master_readdatavalid -> hdd1:sd_master_readdatavalid
	wire         hdd1_avalon_master_write;                                             // hdd1:sd_master_write -> mm_interconnect_1:hdd1_avalon_master_write
	wire  [31:0] hdd1_avalon_master_writedata;                                         // hdd1:sd_master_writedata -> mm_interconnect_1:hdd1_avalon_master_writedata
	wire         mm_bridge_m0_waitrequest;                                             // mm_interconnect_1:mm_bridge_m0_waitrequest -> mm_bridge:m0_waitrequest
	wire  [31:0] mm_bridge_m0_readdata;                                                // mm_interconnect_1:mm_bridge_m0_readdata -> mm_bridge:m0_readdata
	wire         mm_bridge_m0_debugaccess;                                             // mm_bridge:m0_debugaccess -> mm_interconnect_1:mm_bridge_m0_debugaccess
	wire  [31:0] mm_bridge_m0_address;                                                 // mm_bridge:m0_address -> mm_interconnect_1:mm_bridge_m0_address
	wire         mm_bridge_m0_read;                                                    // mm_bridge:m0_read -> mm_interconnect_1:mm_bridge_m0_read
	wire   [3:0] mm_bridge_m0_byteenable;                                              // mm_bridge:m0_byteenable -> mm_interconnect_1:mm_bridge_m0_byteenable
	wire         mm_bridge_m0_readdatavalid;                                           // mm_interconnect_1:mm_bridge_m0_readdatavalid -> mm_bridge:m0_readdatavalid
	wire  [31:0] mm_bridge_m0_writedata;                                               // mm_bridge:m0_writedata -> mm_interconnect_1:mm_bridge_m0_writedata
	wire         mm_bridge_m0_write;                                                   // mm_bridge:m0_write -> mm_interconnect_1:mm_bridge_m0_write
	wire   [0:0] mm_bridge_m0_burstcount;                                              // mm_bridge:m0_burstcount -> mm_interconnect_1:mm_bridge_m0_burstcount
	wire         pc_dma_avalon_master_waitrequest;                                     // mm_interconnect_1:pc_dma_avalon_master_waitrequest -> pc_dma:avm_waitrequest
	wire   [7:0] pc_dma_avalon_master_readdata;                                        // mm_interconnect_1:pc_dma_avalon_master_readdata -> pc_dma:avm_readdata
	wire  [31:0] pc_dma_avalon_master_address;                                         // pc_dma:avm_address -> mm_interconnect_1:pc_dma_avalon_master_address
	wire         pc_dma_avalon_master_read;                                            // pc_dma:avm_read -> mm_interconnect_1:pc_dma_avalon_master_read
	wire         pc_dma_avalon_master_readdatavalid;                                   // mm_interconnect_1:pc_dma_avalon_master_readdatavalid -> pc_dma:avm_readdatavalid
	wire         pc_dma_avalon_master_write;                                           // pc_dma:avm_write -> mm_interconnect_1:pc_dma_avalon_master_write
	wire   [7:0] pc_dma_avalon_master_writedata;                                       // pc_dma:avm_writedata -> mm_interconnect_1:pc_dma_avalon_master_writedata
	wire  [31:0] pc_bus_avalon_sdram_master_readdata;                                  // mm_interconnect_1:pc_bus_avalon_sdram_master_readdata -> pc_bus:sdram_readdata
	wire         pc_bus_avalon_sdram_master_waitrequest;                               // mm_interconnect_1:pc_bus_avalon_sdram_master_waitrequest -> pc_bus:sdram_waitrequest
	wire  [31:0] pc_bus_avalon_sdram_master_address;                                   // pc_bus:sdram_address -> mm_interconnect_1:pc_bus_avalon_sdram_master_address
	wire   [3:0] pc_bus_avalon_sdram_master_byteenable;                                // pc_bus:sdram_byteenable -> mm_interconnect_1:pc_bus_avalon_sdram_master_byteenable
	wire         pc_bus_avalon_sdram_master_read;                                      // pc_bus:sdram_read -> mm_interconnect_1:pc_bus_avalon_sdram_master_read
	wire         pc_bus_avalon_sdram_master_readdatavalid;                             // mm_interconnect_1:pc_bus_avalon_sdram_master_readdatavalid -> pc_bus:sdram_readdatavalid
	wire         pc_bus_avalon_sdram_master_write;                                     // pc_bus:sdram_write -> mm_interconnect_1:pc_bus_avalon_sdram_master_write
	wire  [31:0] pc_bus_avalon_sdram_master_writedata;                                 // pc_bus:sdram_writedata -> mm_interconnect_1:pc_bus_avalon_sdram_master_writedata
	wire   [2:0] pc_bus_avalon_sdram_master_burstcount;                                // pc_bus:sdram_burstcount -> mm_interconnect_1:pc_bus_avalon_sdram_master_burstcount
	wire  [31:0] mm_interconnect_1_driver_sd_avalon_slave_0_readdata;                  // driver_sd:avs_readdata -> mm_interconnect_1:driver_sd_avalon_slave_0_readdata
	wire   [2:0] mm_interconnect_1_driver_sd_avalon_slave_0_address;                   // mm_interconnect_1:driver_sd_avalon_slave_0_address -> driver_sd:avs_address
	wire         mm_interconnect_1_driver_sd_avalon_slave_0_read;                      // mm_interconnect_1:driver_sd_avalon_slave_0_read -> driver_sd:avs_read
	wire         mm_interconnect_1_driver_sd_avalon_slave_0_write;                     // mm_interconnect_1:driver_sd_avalon_slave_0_write -> driver_sd:avs_write
	wire  [31:0] mm_interconnect_1_driver_sd_avalon_slave_0_writedata;                 // mm_interconnect_1:driver_sd_avalon_slave_0_writedata -> driver_sd:avs_writedata
	wire   [1:0] mm_interconnect_1_pc_bus_ctrl_address;                                // mm_interconnect_1:pc_bus_ctrl_address -> pc_bus:ctrl_address
	wire         mm_interconnect_1_pc_bus_ctrl_write;                                  // mm_interconnect_1:pc_bus_ctrl_write -> pc_bus:ctrl_write
	wire  [31:0] mm_interconnect_1_pc_bus_ctrl_writedata;                              // mm_interconnect_1:pc_bus_ctrl_writedata -> pc_bus:ctrl_writedata
	wire   [3:0] mm_interconnect_1_floppy0_mgmt_address;                               // mm_interconnect_1:floppy0_mgmt_address -> floppy0:mgmt_address
	wire         mm_interconnect_1_floppy0_mgmt_write;                                 // mm_interconnect_1:floppy0_mgmt_write -> floppy0:mgmt_write
	wire  [31:0] mm_interconnect_1_floppy0_mgmt_writedata;                             // mm_interconnect_1:floppy0_mgmt_writedata -> floppy0:mgmt_writedata
	wire   [2:0] mm_interconnect_1_hdd0_mgmt_address;                                  // mm_interconnect_1:hdd0_mgmt_address -> hdd0:mgmt_address
	wire         mm_interconnect_1_hdd0_mgmt_write;                                    // mm_interconnect_1:hdd0_mgmt_write -> hdd0:mgmt_write
	wire  [31:0] mm_interconnect_1_hdd0_mgmt_writedata;                                // mm_interconnect_1:hdd0_mgmt_writedata -> hdd0:mgmt_writedata
	wire   [7:0] mm_interconnect_1_rtc_mgmt_address;                                   // mm_interconnect_1:rtc_mgmt_address -> rtc:mgmt_address
	wire         mm_interconnect_1_rtc_mgmt_write;                                     // mm_interconnect_1:rtc_mgmt_write -> rtc:mgmt_write
	wire  [31:0] mm_interconnect_1_rtc_mgmt_writedata;                                 // mm_interconnect_1:rtc_mgmt_writedata -> rtc:mgmt_writedata
	wire   [8:0] mm_interconnect_1_sound_mgmt_address;                                 // mm_interconnect_1:sound_mgmt_address -> sound:mgmt_address
	wire         mm_interconnect_1_sound_mgmt_write;                                   // mm_interconnect_1:sound_mgmt_write -> sound:mgmt_write
	wire  [31:0] mm_interconnect_1_sound_mgmt_writedata;                               // mm_interconnect_1:sound_mgmt_writedata -> sound:mgmt_writedata
	wire   [0:0] mm_interconnect_1_pit_mgmt_address;                                   // mm_interconnect_1:pit_mgmt_address -> pit:mgmt_address
	wire         mm_interconnect_1_pit_mgmt_write;                                     // mm_interconnect_1:pit_mgmt_write -> pit:mgmt_write
	wire  [31:0] mm_interconnect_1_pit_mgmt_writedata;                                 // mm_interconnect_1:pit_mgmt_writedata -> pit:mgmt_writedata
	wire   [2:0] mm_interconnect_1_hdd1_mgmt_address;                                  // mm_interconnect_1:hdd1_mgmt_address -> hdd1:mgmt_address
	wire         mm_interconnect_1_hdd1_mgmt_write;                                    // mm_interconnect_1:hdd1_mgmt_write -> hdd1:mgmt_write
	wire  [31:0] mm_interconnect_1_hdd1_mgmt_writedata;                                // mm_interconnect_1:hdd1_mgmt_writedata -> hdd1:mgmt_writedata
	wire   [7:0] mm_interconnect_1_floppy0_sd_slave_readdata;                          // floppy0:sd_slave_readdata -> mm_interconnect_1:floppy0_sd_slave_readdata
	wire   [8:0] mm_interconnect_1_floppy0_sd_slave_address;                           // mm_interconnect_1:floppy0_sd_slave_address -> floppy0:sd_slave_address
	wire         mm_interconnect_1_floppy0_sd_slave_read;                              // mm_interconnect_1:floppy0_sd_slave_read -> floppy0:sd_slave_read
	wire         mm_interconnect_1_floppy0_sd_slave_write;                             // mm_interconnect_1:floppy0_sd_slave_write -> floppy0:sd_slave_write
	wire   [7:0] mm_interconnect_1_floppy0_sd_slave_writedata;                         // mm_interconnect_1:floppy0_sd_slave_writedata -> floppy0:sd_slave_writedata
	wire  [31:0] mm_interconnect_1_hdd0_sd_slave_readdata;                             // hdd0:sd_slave_readdata -> mm_interconnect_1:hdd0_sd_slave_readdata
	wire   [8:0] mm_interconnect_1_hdd0_sd_slave_address;                              // mm_interconnect_1:hdd0_sd_slave_address -> hdd0:sd_slave_address
	wire         mm_interconnect_1_hdd0_sd_slave_read;                                 // mm_interconnect_1:hdd0_sd_slave_read -> hdd0:sd_slave_read
	wire         mm_interconnect_1_hdd0_sd_slave_write;                                // mm_interconnect_1:hdd0_sd_slave_write -> hdd0:sd_slave_write
	wire  [31:0] mm_interconnect_1_hdd0_sd_slave_writedata;                            // mm_interconnect_1:hdd0_sd_slave_writedata -> hdd0:sd_slave_writedata
	wire  [31:0] mm_interconnect_1_hdd1_sd_slave_readdata;                             // hdd1:sd_slave_readdata -> mm_interconnect_1:hdd1_sd_slave_readdata
	wire   [8:0] mm_interconnect_1_hdd1_sd_slave_address;                              // mm_interconnect_1:hdd1_sd_slave_address -> hdd1:sd_slave_address
	wire         mm_interconnect_1_hdd1_sd_slave_read;                                 // mm_interconnect_1:hdd1_sd_slave_read -> hdd1:sd_slave_read
	wire         mm_interconnect_1_hdd1_sd_slave_write;                                // mm_interconnect_1:hdd1_sd_slave_write -> hdd1:sd_slave_write
	wire  [31:0] mm_interconnect_1_hdd1_sd_slave_writedata;                            // mm_interconnect_1:hdd1_sd_slave_writedata -> hdd1:sd_slave_writedata
	wire  [63:0] mm_interconnect_1_address_span_extender_windowed_slave_readdata;      // address_span_extender:avs_s0_readdata -> mm_interconnect_1:address_span_extender_windowed_slave_readdata
	wire         mm_interconnect_1_address_span_extender_windowed_slave_waitrequest;   // address_span_extender:avs_s0_waitrequest -> mm_interconnect_1:address_span_extender_windowed_slave_waitrequest
	wire  [23:0] mm_interconnect_1_address_span_extender_windowed_slave_address;       // mm_interconnect_1:address_span_extender_windowed_slave_address -> address_span_extender:avs_s0_address
	wire         mm_interconnect_1_address_span_extender_windowed_slave_read;          // mm_interconnect_1:address_span_extender_windowed_slave_read -> address_span_extender:avs_s0_read
	wire   [7:0] mm_interconnect_1_address_span_extender_windowed_slave_byteenable;    // mm_interconnect_1:address_span_extender_windowed_slave_byteenable -> address_span_extender:avs_s0_byteenable
	wire         mm_interconnect_1_address_span_extender_windowed_slave_readdatavalid; // address_span_extender:avs_s0_readdatavalid -> mm_interconnect_1:address_span_extender_windowed_slave_readdatavalid
	wire         mm_interconnect_1_address_span_extender_windowed_slave_write;         // mm_interconnect_1:address_span_extender_windowed_slave_write -> address_span_extender:avs_s0_write
	wire  [63:0] mm_interconnect_1_address_span_extender_windowed_slave_writedata;     // mm_interconnect_1:address_span_extender_windowed_slave_writedata -> address_span_extender:avs_s0_writedata
	wire   [7:0] mm_interconnect_1_address_span_extender_windowed_slave_burstcount;    // mm_interconnect_1:address_span_extender_windowed_slave_burstcount -> address_span_extender:avs_s0_burstcount
	wire  [31:0] pc_bus_avalon_vga_master_readdata;                                    // mm_interconnect_3:pc_bus_avalon_vga_master_readdata -> pc_bus:vga_readdata
	wire         pc_bus_avalon_vga_master_waitrequest;                                 // mm_interconnect_3:pc_bus_avalon_vga_master_waitrequest -> pc_bus:vga_waitrequest
	wire  [31:0] pc_bus_avalon_vga_master_address;                                     // pc_bus:vga_address -> mm_interconnect_3:pc_bus_avalon_vga_master_address
	wire   [3:0] pc_bus_avalon_vga_master_byteenable;                                  // pc_bus:vga_byteenable -> mm_interconnect_3:pc_bus_avalon_vga_master_byteenable
	wire         pc_bus_avalon_vga_master_read;                                        // pc_bus:vga_read -> mm_interconnect_3:pc_bus_avalon_vga_master_read
	wire         pc_bus_avalon_vga_master_readdatavalid;                               // mm_interconnect_3:pc_bus_avalon_vga_master_readdatavalid -> pc_bus:vga_readdatavalid
	wire         pc_bus_avalon_vga_master_write;                                       // pc_bus:vga_write -> mm_interconnect_3:pc_bus_avalon_vga_master_write
	wire  [31:0] pc_bus_avalon_vga_master_writedata;                                   // pc_bus:vga_writedata -> mm_interconnect_3:pc_bus_avalon_vga_master_writedata
	wire   [2:0] pc_bus_avalon_vga_master_burstcount;                                  // pc_bus:vga_burstcount -> mm_interconnect_3:pc_bus_avalon_vga_master_burstcount
	wire   [7:0] mm_interconnect_3_vga_mem_readdata;                                   // vga:mem_readdata -> mm_interconnect_3:vga_mem_readdata
	wire  [16:0] mm_interconnect_3_vga_mem_address;                                    // mm_interconnect_3:vga_mem_address -> vga:mem_address
	wire         mm_interconnect_3_vga_mem_read;                                       // mm_interconnect_3:vga_mem_read -> vga:mem_read
	wire         mm_interconnect_3_vga_mem_write;                                      // mm_interconnect_3:vga_mem_write -> vga:mem_write
	wire   [7:0] mm_interconnect_3_vga_mem_writedata;                                  // mm_interconnect_3:vga_mem_writedata -> vga:mem_writedata
	wire         irq_mapper_receiver0_irq;                                             // pit:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                             // rtc:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                             // sound:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                             // hdd0:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                             // floppy0:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                             // hdd1:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                             // vga:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                             // ps2:irq_keyb -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                             // ps2:irq_mouse -> irq_mapper:receiver8_irq
	wire  [15:0] pic_interrupt_receiver_irq;                                           // irq_mapper:sender_irq -> pic:interrupt_input
	wire         irq_mapper_receiver9_irq;                                             // irq_synchronizer:sender_irq -> irq_mapper:receiver9_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                        // uart:intr -> irq_synchronizer:receiver_irq
	wire         rst_controller_reset_out_reset;                                       // rst_controller:reset_out -> [ao486:rst_n, mm_interconnect_0:ao486_reset_sink_reset_bridge_in_reset_reset]
	wire         rst_controller_001_reset_out_reset;                                   // rst_controller_001:reset_out -> [irq_synchronizer:receiver_reset, mm_interconnect_0:width_trans_reset_reset_bridge_in_reset_reset, uart:rst_n, width_trans:reset]

	altera_address_span_extender #(
		.DATA_WIDTH           (64),
		.BYTEENABLE_WIDTH     (8),
		.MASTER_ADDRESS_WIDTH (32),
		.SLAVE_ADDRESS_WIDTH  (24),
		.SLAVE_ADDRESS_SHIFT  (3),
		.BURSTCOUNT_WIDTH     (8),
		.CNTL_ADDRESS_WIDTH   (1),
		.SUB_WINDOW_COUNT     (1),
		.MASTER_ADDRESS_DEF   (64'b0000000000000000000000000000000000110000000000000000000000000000)
	) address_span_extender (
		.clk                  (clk_sys_clk),                                                          //           clock.clk
		.reset                (reset_sys_reset_out_reset),                                            //           reset.reset
		.avs_s0_address       (mm_interconnect_1_address_span_extender_windowed_slave_address),       //  windowed_slave.address
		.avs_s0_read          (mm_interconnect_1_address_span_extender_windowed_slave_read),          //                .read
		.avs_s0_readdata      (mm_interconnect_1_address_span_extender_windowed_slave_readdata),      //                .readdata
		.avs_s0_write         (mm_interconnect_1_address_span_extender_windowed_slave_write),         //                .write
		.avs_s0_writedata     (mm_interconnect_1_address_span_extender_windowed_slave_writedata),     //                .writedata
		.avs_s0_readdatavalid (mm_interconnect_1_address_span_extender_windowed_slave_readdatavalid), //                .readdatavalid
		.avs_s0_waitrequest   (mm_interconnect_1_address_span_extender_windowed_slave_waitrequest),   //                .waitrequest
		.avs_s0_byteenable    (mm_interconnect_1_address_span_extender_windowed_slave_byteenable),    //                .byteenable
		.avs_s0_burstcount    (mm_interconnect_1_address_span_extender_windowed_slave_burstcount),    //                .burstcount
		.avm_m0_address       (ddram_address),                                                        // expanded_master.address
		.avm_m0_read          (ddram_read),                                                           //                .read
		.avm_m0_waitrequest   (ddram_waitrequest),                                                    //                .waitrequest
		.avm_m0_readdata      (ddram_readdata),                                                       //                .readdata
		.avm_m0_write         (ddram_write),                                                          //                .write
		.avm_m0_writedata     (ddram_writedata),                                                      //                .writedata
		.avm_m0_readdatavalid (ddram_readdatavalid),                                                  //                .readdatavalid
		.avm_m0_byteenable    (ddram_byteenable),                                                     //                .byteenable
		.avm_m0_burstcount    (ddram_burstcount),                                                     //                .burstcount
		.avs_cntl_address     (1'b0),                                                                 //     (terminated)
		.avs_cntl_read        (1'b0),                                                                 //     (terminated)
		.avs_cntl_readdata    (),                                                                     //     (terminated)
		.avs_cntl_write       (1'b0),                                                                 //     (terminated)
		.avs_cntl_writedata   (64'b0000000000000000000000000000000000000000000000000000000000000000), //     (terminated)
		.avs_cntl_byteenable  (8'b00000000)                                                           //     (terminated)
	);

	ao486 ao486 (
		.clk                     (clk_sys_clk),                            //         clock.clk
		.rst_n                   (~rst_controller_reset_out_reset),        //    reset_sink.reset_n
		.avm_address             (ao486_avalon_memory_address),            // avalon_memory.address
		.avm_writedata           (ao486_avalon_memory_writedata),          //              .writedata
		.avm_byteenable          (ao486_avalon_memory_byteenable),         //              .byteenable
		.avm_burstcount          (ao486_avalon_memory_burstcount),         //              .burstcount
		.avm_write               (ao486_avalon_memory_write),              //              .write
		.avm_read                (ao486_avalon_memory_read),               //              .read
		.avm_waitrequest         (ao486_avalon_memory_waitrequest),        //              .waitrequest
		.avm_readdatavalid       (ao486_avalon_memory_readdatavalid),      //              .readdatavalid
		.avm_readdata            (ao486_avalon_memory_readdata),           //              .readdata
		.interrupt_do            (pic_conduit_interrupt_interrupt_do),     //     interrupt.interrupt_do
		.interrupt_vector        (pic_conduit_interrupt_interrupt_vector), //              .interrupt_vector
		.interrupt_done          (ao486_interrupt_interrupt_done),         //              .interrupt_done
		.avalon_io_address       (ao486_avalon_io_address),                //     avalon_io.address
		.avalon_io_byteenable    (ao486_avalon_io_byteenable),             //              .byteenable
		.avalon_io_read          (ao486_avalon_io_read),                   //              .read
		.avalon_io_readdatavalid (ao486_avalon_io_readdatavalid),          //              .readdatavalid
		.avalon_io_readdata      (ao486_avalon_io_readdata),               //              .readdata
		.avalon_io_write         (ao486_avalon_io_write),                  //              .write
		.avalon_io_writedata     (ao486_avalon_io_writedata),              //              .writedata
		.avalon_io_waitrequest   (ao486_avalon_io_waitrequest),            //              .waitrequest
		.a20_enable              (ps2_conduit_a20_a20_enable)              //   conduit_a20.a20_enable
	);

	driver_sd driver_sd (
		.clk           (clk_sys_clk),                                          //          clock.clk
		.avs_address   (mm_interconnect_1_driver_sd_avalon_slave_0_address),   // avalon_slave_0.address
		.avs_read      (mm_interconnect_1_driver_sd_avalon_slave_0_read),      //               .read
		.avs_readdata  (mm_interconnect_1_driver_sd_avalon_slave_0_readdata),  //               .readdata
		.avs_write     (mm_interconnect_1_driver_sd_avalon_slave_0_write),     //               .write
		.avs_writedata (mm_interconnect_1_driver_sd_avalon_slave_0_writedata), //               .writedata
		.rst_n         (~reset_sys_reset_out_reset),                           //     reset_sink.reset_n
		.op_read       (disk_op_read),                                         //    conduit_prx.op_read
		.op_write      (disk_op_write),                                        //               .op_write
		.result_ok     (disk_result_ok),                                       //               .result_ok
		.result_error  (disk_result_error),                                    //               .result_error
		.op_device     (disk_op_device)                                        //               .op_device
	);

	floppy #(
		.BufAddress (32'b00000000000000000000100000000000)
	) floppy0 (
		.clk                     (clk_sys_clk),                                     //              clock.clk
		.io_address              (mm_interconnect_0_floppy0_io_address),            //                 io.address
		.io_read                 (mm_interconnect_0_floppy0_io_read),               //                   .read
		.io_readdata             (mm_interconnect_0_floppy0_io_readdata),           //                   .readdata
		.io_write                (mm_interconnect_0_floppy0_io_write),              //                   .write
		.io_writedata            (mm_interconnect_0_floppy0_io_writedata),          //                   .writedata
		.sd_slave_address        (mm_interconnect_1_floppy0_sd_slave_address),      //           sd_slave.address
		.sd_slave_read           (mm_interconnect_1_floppy0_sd_slave_read),         //                   .read
		.sd_slave_readdata       (mm_interconnect_1_floppy0_sd_slave_readdata),     //                   .readdata
		.sd_slave_write          (mm_interconnect_1_floppy0_sd_slave_write),        //                   .write
		.sd_slave_writedata      (mm_interconnect_1_floppy0_sd_slave_writedata),    //                   .writedata
		.mgmt_address            (mm_interconnect_1_floppy0_mgmt_address),          //               mgmt.address
		.mgmt_write              (mm_interconnect_1_floppy0_mgmt_write),            //                   .write
		.mgmt_writedata          (mm_interconnect_1_floppy0_mgmt_writedata),        //                   .writedata
		.rst_n                   (~reset_sys_reset_out_reset),                      //         reset_sink.reset_n
		.sd_master_address       (floppy0_avalon_master_address),                   //      avalon_master.address
		.sd_master_waitrequest   (floppy0_avalon_master_waitrequest),               //                   .waitrequest
		.sd_master_read          (floppy0_avalon_master_read),                      //                   .read
		.sd_master_readdatavalid (floppy0_avalon_master_readdatavalid),             //                   .readdatavalid
		.sd_master_readdata      (floppy0_avalon_master_readdata),                  //                   .readdata
		.sd_master_write         (floppy0_avalon_master_write),                     //                   .write
		.sd_master_writedata     (floppy0_avalon_master_writedata),                 //                   .writedata
		.dma_floppy_req          (floppy0_conduit_dma_floppy_dma_floppy_req),       // conduit_dma_floppy.dma_floppy_req
		.dma_floppy_ack          (pc_dma_conduit_dma_floppy_dma_floppy_ack),        //                   .dma_floppy_ack
		.dma_floppy_terminal     (pc_dma_conduit_dma_floppy_dma_floppy_terminal),   //                   .dma_floppy_terminal
		.dma_floppy_readdata     (pc_dma_conduit_dma_floppy_dma_floppy_readdata),   //                   .dma_floppy_readdata
		.dma_floppy_writedata    (floppy0_conduit_dma_floppy_dma_floppy_writedata), //                   .dma_floppy_writedata
		.ide_3f6_read            (floppy0_conduit_ide_3f6_ide_3f6_read),            //    conduit_ide_3f6.ide_3f6_read
		.ide_3f6_readdata        (hdd0_conduit_ide_3f6_ide_3f6_readdata),           //                   .ide_3f6_readdata
		.ide_3f6_write           (floppy0_conduit_ide_3f6_ide_3f6_write),           //                   .ide_3f6_write
		.ide_3f6_writedata       (floppy0_conduit_ide_3f6_ide_3f6_writedata),       //                   .ide_3f6_writedata
		.irq                     (irq_mapper_receiver4_irq)                         //   interrupt_sender.irq
	);

	hdd #(
		.BufAddress (32'b00000000000000000000000000000000)
	) hdd0 (
		.clk                     (clk_sys_clk),                               //            clock.clk
		.io_address              (mm_interconnect_0_hdd0_io_address),         //               io.address
		.io_byteenable           (mm_interconnect_0_hdd0_io_byteenable),      //                 .byteenable
		.io_read                 (mm_interconnect_0_hdd0_io_read),            //                 .read
		.io_readdata             (mm_interconnect_0_hdd0_io_readdata),        //                 .readdata
		.io_write                (mm_interconnect_0_hdd0_io_write),           //                 .write
		.io_writedata            (mm_interconnect_0_hdd0_io_writedata),       //                 .writedata
		.sd_slave_address        (mm_interconnect_1_hdd0_sd_slave_address),   //         sd_slave.address
		.sd_slave_read           (mm_interconnect_1_hdd0_sd_slave_read),      //                 .read
		.sd_slave_readdata       (mm_interconnect_1_hdd0_sd_slave_readdata),  //                 .readdata
		.sd_slave_write          (mm_interconnect_1_hdd0_sd_slave_write),     //                 .write
		.sd_slave_writedata      (mm_interconnect_1_hdd0_sd_slave_writedata), //                 .writedata
		.mgmt_address            (mm_interconnect_1_hdd0_mgmt_address),       //             mgmt.address
		.mgmt_write              (mm_interconnect_1_hdd0_mgmt_write),         //                 .write
		.mgmt_writedata          (mm_interconnect_1_hdd0_mgmt_writedata),     //                 .writedata
		.rst_n                   (~reset_sys_reset_out_reset),                //       reset_sink.reset_n
		.irq                     (irq_mapper_receiver3_irq),                  // interrupt_sender.irq
		.sd_master_address       (hdd0_avalon_master_address),                //    avalon_master.address
		.sd_master_waitrequest   (hdd0_avalon_master_waitrequest),            //                 .waitrequest
		.sd_master_read          (hdd0_avalon_master_read),                   //                 .read
		.sd_master_readdatavalid (hdd0_avalon_master_readdatavalid),          //                 .readdatavalid
		.sd_master_readdata      (hdd0_avalon_master_readdata),               //                 .readdata
		.sd_master_write         (hdd0_avalon_master_write),                  //                 .write
		.sd_master_writedata     (hdd0_avalon_master_writedata),              //                 .writedata
		.ide_3f6_read            (floppy0_conduit_ide_3f6_ide_3f6_read),      //  conduit_ide_3f6.ide_3f6_read
		.ide_3f6_readdata        (hdd0_conduit_ide_3f6_ide_3f6_readdata),     //                 .ide_3f6_readdata
		.ide_3f6_write           (floppy0_conduit_ide_3f6_ide_3f6_write),     //                 .ide_3f6_write
		.ide_3f6_writedata       (floppy0_conduit_ide_3f6_ide_3f6_writedata)  //                 .ide_3f6_writedata
	);

	hdd #(
		.BufAddress (32'b00000000000000000001000000000000)
	) hdd1 (
		.clk                     (clk_sys_clk),                                    //            clock.clk
		.io_address              (mm_interconnect_0_hdd1_io_address),              //               io.address
		.io_byteenable           (mm_interconnect_0_hdd1_io_byteenable),           //                 .byteenable
		.io_read                 (mm_interconnect_0_hdd1_io_read),                 //                 .read
		.io_readdata             (mm_interconnect_0_hdd1_io_readdata),             //                 .readdata
		.io_write                (mm_interconnect_0_hdd1_io_write),                //                 .write
		.io_writedata            (mm_interconnect_0_hdd1_io_writedata),            //                 .writedata
		.sd_slave_address        (mm_interconnect_1_hdd1_sd_slave_address),        //         sd_slave.address
		.sd_slave_read           (mm_interconnect_1_hdd1_sd_slave_read),           //                 .read
		.sd_slave_readdata       (mm_interconnect_1_hdd1_sd_slave_readdata),       //                 .readdata
		.sd_slave_write          (mm_interconnect_1_hdd1_sd_slave_write),          //                 .write
		.sd_slave_writedata      (mm_interconnect_1_hdd1_sd_slave_writedata),      //                 .writedata
		.mgmt_address            (mm_interconnect_1_hdd1_mgmt_address),            //             mgmt.address
		.mgmt_write              (mm_interconnect_1_hdd1_mgmt_write),              //                 .write
		.mgmt_writedata          (mm_interconnect_1_hdd1_mgmt_writedata),          //                 .writedata
		.rst_n                   (~reset_sys_reset_out_reset),                     //       reset_sink.reset_n
		.irq                     (irq_mapper_receiver5_irq),                       // interrupt_sender.irq
		.sd_master_address       (hdd1_avalon_master_address),                     //    avalon_master.address
		.sd_master_waitrequest   (hdd1_avalon_master_waitrequest),                 //                 .waitrequest
		.sd_master_read          (hdd1_avalon_master_read),                        //                 .read
		.sd_master_readdatavalid (hdd1_avalon_master_readdatavalid),               //                 .readdatavalid
		.sd_master_readdata      (hdd1_avalon_master_readdata),                    //                 .readdata
		.sd_master_write         (hdd1_avalon_master_write),                       //                 .write
		.sd_master_writedata     (hdd1_avalon_master_writedata),                   //                 .writedata
		.ide_3f6_read            (hddext_0x370_conduit_ide_3f6_ide_3f6_read),      //  conduit_ide_3f6.ide_3f6_read
		.ide_3f6_readdata        (hdd1_conduit_ide_3f6_ide_3f6_readdata),          //                 .ide_3f6_readdata
		.ide_3f6_write           (hddext_0x370_conduit_ide_3f6_ide_3f6_write),     //                 .ide_3f6_write
		.ide_3f6_writedata       (hddext_0x370_conduit_ide_3f6_ide_3f6_writedata)  //                 .ide_3f6_writedata
	);

	hddext hddext_0x370 (
		.clk               (clk_sys_clk),                                    //           clock.clk
		.io_address        (mm_interconnect_0_hddext_0x370_io_address),      //              io.address
		.io_read           (mm_interconnect_0_hddext_0x370_io_read),         //                .read
		.io_readdata       (mm_interconnect_0_hddext_0x370_io_readdata),     //                .readdata
		.io_write          (mm_interconnect_0_hddext_0x370_io_write),        //                .write
		.io_writedata      (mm_interconnect_0_hddext_0x370_io_writedata),    //                .writedata
		.rst_n             (~reset_sys_reset_out_reset),                     //      reset_sink.reset_n
		.ide_3f6_read      (hddext_0x370_conduit_ide_3f6_ide_3f6_read),      // conduit_ide_3f6.ide_3f6_read
		.ide_3f6_readdata  (hdd1_conduit_ide_3f6_ide_3f6_readdata),          //                .ide_3f6_readdata
		.ide_3f6_write     (hddext_0x370_conduit_ide_3f6_ide_3f6_write),     //                .ide_3f6_write
		.ide_3f6_writedata (hddext_0x370_conduit_ide_3f6_ide_3f6_writedata)  //                .ide_3f6_writedata
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (32),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) mm_bridge (
		.clk              (clk_sys_clk),                //   clk.clk
		.reset            (reset_sys_reset_out_reset),  // reset.reset
		.s0_waitrequest   (mem_waitrequest),            //    s0.waitrequest
		.s0_readdata      (mem_readdata),               //      .readdata
		.s0_readdatavalid (mem_readdatavalid),          //      .readdatavalid
		.s0_burstcount    (mem_burstcount),             //      .burstcount
		.s0_writedata     (mem_writedata),              //      .writedata
		.s0_address       (mem_address),                //      .address
		.s0_write         (mem_write),                  //      .write
		.s0_read          (mem_read),                   //      .read
		.s0_byteenable    (mem_byteenable),             //      .byteenable
		.s0_debugaccess   (mem_debugaccess),            //      .debugaccess
		.m0_waitrequest   (mm_bridge_m0_waitrequest),   //    m0.waitrequest
		.m0_readdata      (mm_bridge_m0_readdata),      //      .readdata
		.m0_readdatavalid (mm_bridge_m0_readdatavalid), //      .readdatavalid
		.m0_burstcount    (mm_bridge_m0_burstcount),    //      .burstcount
		.m0_writedata     (mm_bridge_m0_writedata),     //      .writedata
		.m0_address       (mm_bridge_m0_address),       //      .address
		.m0_write         (mm_bridge_m0_write),         //      .write
		.m0_read          (mm_bridge_m0_read),          //      .read
		.m0_byteenable    (mm_bridge_m0_byteenable),    //      .byteenable
		.m0_debugaccess   (mm_bridge_m0_debugaccess),   //      .debugaccess
		.s0_response      (),                           // (terminated)
		.m0_response      (2'b00)                       // (terminated)
	);

	pc_bus pc_bus (
		.clk                 (clk_sys_clk),                              //               clock.clk
		.ctrl_address        (mm_interconnect_1_pc_bus_ctrl_address),    //                ctrl.address
		.ctrl_write          (mm_interconnect_1_pc_bus_ctrl_write),      //                    .write
		.ctrl_writedata      (mm_interconnect_1_pc_bus_ctrl_writedata),  //                    .writedata
		.mem_address         (ao486_avalon_memory_address),              //                 mem.address
		.mem_byteenable      (ao486_avalon_memory_byteenable),           //                    .byteenable
		.mem_read            (ao486_avalon_memory_read),                 //                    .read
		.mem_readdata        (ao486_avalon_memory_readdata),             //                    .readdata
		.mem_write           (ao486_avalon_memory_write),                //                    .write
		.mem_writedata       (ao486_avalon_memory_writedata),            //                    .writedata
		.mem_waitrequest     (ao486_avalon_memory_waitrequest),          //                    .waitrequest
		.mem_readdatavalid   (ao486_avalon_memory_readdatavalid),        //                    .readdatavalid
		.mem_burstcount      (ao486_avalon_memory_burstcount),           //                    .burstcount
		.rst_n               (~reset_sys_reset_out_reset),               //          reset_sink.reset_n
		.vga_address         (pc_bus_avalon_vga_master_address),         //   avalon_vga_master.address
		.vga_byteenable      (pc_bus_avalon_vga_master_byteenable),      //                    .byteenable
		.vga_read            (pc_bus_avalon_vga_master_read),            //                    .read
		.vga_readdata        (pc_bus_avalon_vga_master_readdata),        //                    .readdata
		.vga_write           (pc_bus_avalon_vga_master_write),           //                    .write
		.vga_writedata       (pc_bus_avalon_vga_master_writedata),       //                    .writedata
		.vga_waitrequest     (pc_bus_avalon_vga_master_waitrequest),     //                    .waitrequest
		.vga_readdatavalid   (pc_bus_avalon_vga_master_readdatavalid),   //                    .readdatavalid
		.vga_burstcount      (pc_bus_avalon_vga_master_burstcount),      //                    .burstcount
		.sdram_address       (pc_bus_avalon_sdram_master_address),       // avalon_sdram_master.address
		.sdram_byteenable    (pc_bus_avalon_sdram_master_byteenable),    //                    .byteenable
		.sdram_read          (pc_bus_avalon_sdram_master_read),          //                    .read
		.sdram_readdata      (pc_bus_avalon_sdram_master_readdata),      //                    .readdata
		.sdram_write         (pc_bus_avalon_sdram_master_write),         //                    .write
		.sdram_writedata     (pc_bus_avalon_sdram_master_writedata),     //                    .writedata
		.sdram_waitrequest   (pc_bus_avalon_sdram_master_waitrequest),   //                    .waitrequest
		.sdram_readdatavalid (pc_bus_avalon_sdram_master_readdatavalid), //                    .readdatavalid
		.sdram_burstcount    (pc_bus_avalon_sdram_master_burstcount)     //                    .burstcount
	);

	pc_dma pc_dma (
		.clk                        (clk_sys_clk),                                               //                    clock.clk
		.slave_address              (mm_interconnect_0_pc_dma_slave_address),                    //                    slave.address
		.slave_read                 (mm_interconnect_0_pc_dma_slave_read),                       //                         .read
		.slave_readdata             (mm_interconnect_0_pc_dma_slave_readdata),                   //                         .readdata
		.slave_write                (mm_interconnect_0_pc_dma_slave_write),                      //                         .write
		.slave_writedata            (mm_interconnect_0_pc_dma_slave_writedata),                  //                         .writedata
		.page_address               (mm_interconnect_0_pc_dma_page_address),                     //                     page.address
		.page_read                  (mm_interconnect_0_pc_dma_page_read),                        //                         .read
		.page_readdata              (mm_interconnect_0_pc_dma_page_readdata),                    //                         .readdata
		.page_write                 (mm_interconnect_0_pc_dma_page_write),                       //                         .write
		.page_writedata             (mm_interconnect_0_pc_dma_page_writedata),                   //                         .writedata
		.master_address             (mm_interconnect_0_pc_dma_master_address),                   //                   master.address
		.master_read                (mm_interconnect_0_pc_dma_master_read),                      //                         .read
		.master_readdata            (mm_interconnect_0_pc_dma_master_readdata),                  //                         .readdata
		.master_write               (mm_interconnect_0_pc_dma_master_write),                     //                         .write
		.master_writedata           (mm_interconnect_0_pc_dma_master_writedata),                 //                         .writedata
		.rst_n                      (~reset_sys_reset_out_reset),                                //               reset_sink.reset_n
		.avm_address                (pc_dma_avalon_master_address),                              //            avalon_master.address
		.avm_waitrequest            (pc_dma_avalon_master_waitrequest),                          //                         .waitrequest
		.avm_read                   (pc_dma_avalon_master_read),                                 //                         .read
		.avm_readdatavalid          (pc_dma_avalon_master_readdatavalid),                        //                         .readdatavalid
		.avm_readdata               (pc_dma_avalon_master_readdata),                             //                         .readdata
		.avm_write                  (pc_dma_avalon_master_write),                                //                         .write
		.avm_writedata              (pc_dma_avalon_master_writedata),                            //                         .writedata
		.dma_floppy_req             (floppy0_conduit_dma_floppy_dma_floppy_req),                 //       conduit_dma_floppy.dma_floppy_req
		.dma_floppy_ack             (pc_dma_conduit_dma_floppy_dma_floppy_ack),                  //                         .dma_floppy_ack
		.dma_floppy_terminal        (pc_dma_conduit_dma_floppy_dma_floppy_terminal),             //                         .dma_floppy_terminal
		.dma_floppy_readdata        (pc_dma_conduit_dma_floppy_dma_floppy_readdata),             //                         .dma_floppy_readdata
		.dma_floppy_writedata       (floppy0_conduit_dma_floppy_dma_floppy_writedata),           //                         .dma_floppy_writedata
		.dma_soundblaster_req       (sound_conduit_dma_soundblaster_dma_soundblaster_req),       // conduit_dma_soundblaster.dma_soundblaster_req
		.dma_soundblaster_ack       (pc_dma_conduit_dma_soundblaster_dma_soundblaster_ack),      //                         .dma_soundblaster_ack
		.dma_soundblaster_terminal  (pc_dma_conduit_dma_soundblaster_dma_soundblaster_terminal), //                         .dma_soundblaster_terminal
		.dma_soundblaster_readdata  (pc_dma_conduit_dma_soundblaster_dma_soundblaster_readdata), //                         .dma_soundblaster_readdata
		.dma_soundblaster_writedata (sound_conduit_dma_soundblaster_dma_soundblaster_writedata)  //                         .dma_soundblaster_writedata
	);

	pic pic (
		.clk              (clk_sys_clk),                            //              clock.clk
		.master_address   (mm_interconnect_0_pic_master_address),   //             master.address
		.master_read      (mm_interconnect_0_pic_master_read),      //                   .read
		.master_readdata  (mm_interconnect_0_pic_master_readdata),  //                   .readdata
		.master_write     (mm_interconnect_0_pic_master_write),     //                   .write
		.master_writedata (mm_interconnect_0_pic_master_writedata), //                   .writedata
		.slave_address    (mm_interconnect_0_pic_slave_address),    //              slave.address
		.slave_read       (mm_interconnect_0_pic_slave_read),       //                   .read
		.slave_readdata   (mm_interconnect_0_pic_slave_readdata),   //                   .readdata
		.slave_write      (mm_interconnect_0_pic_slave_write),      //                   .write
		.slave_writedata  (mm_interconnect_0_pic_slave_writedata),  //                   .writedata
		.rst_n            (~reset_sys_reset_out_reset),             //         reset_sink.reset_n
		.interrupt_vector (pic_conduit_interrupt_interrupt_vector), //  conduit_interrupt.interrupt_vector
		.interrupt_done   (ao486_interrupt_interrupt_done),         //                   .interrupt_done
		.interrupt_do     (pic_conduit_interrupt_interrupt_do),     //                   .interrupt_do
		.interrupt_input  (pic_interrupt_receiver_irq)              // interrupt_receiver.irq
	);

	pit pit (
		.clk                   (clk_sys_clk),                                   //               clock.clk
		.io_address            (mm_interconnect_0_pit_io_address),              //                  io.address
		.io_read               (mm_interconnect_0_pit_io_read),                 //                    .read
		.io_readdata           (mm_interconnect_0_pit_io_readdata),             //                    .readdata
		.io_write              (mm_interconnect_0_pit_io_write),                //                    .write
		.io_writedata          (mm_interconnect_0_pit_io_writedata),            //                    .writedata
		.mgmt_address          (mm_interconnect_1_pit_mgmt_address),            //                mgmt.address
		.mgmt_write            (mm_interconnect_1_pit_mgmt_write),              //                    .write
		.mgmt_writedata        (mm_interconnect_1_pit_mgmt_writedata),          //                    .writedata
		.rst_n                 (~reset_sys_reset_out_reset),                    //          reset_sink.reset_n
		.speaker_61h_read      (ps2_conduit_speaker_61h_speaker_61h_read),      // conduit_speaker_61h.speaker_61h_read
		.speaker_61h_readdata  (pit_conduit_speaker_61h_speaker_61h_readdata),  //                    .speaker_61h_readdata
		.speaker_61h_write     (ps2_conduit_speaker_61h_speaker_61h_write),     //                    .speaker_61h_write
		.speaker_61h_writedata (ps2_conduit_speaker_61h_speaker_61h_writedata), //                    .speaker_61h_writedata
		.speaker_enable        (speaker_enable),                                //     conduit_speaker.enable
		.speaker_out           (speaker_out),                                   //                    .out
		.irq                   (irq_mapper_receiver0_irq)                       //       interrupt_pit.irq
	);

	system_pll_0 pll_0 (
		.refclk   (clk_clk),           //  refclk.clk
		.rst      (pll_reset_reset),   //   reset.reset
		.outclk_0 (clk_sys_clk),       // outclk0.clk
		.outclk_1 (pll_0_outclk1_clk), // outclk1.clk
		.outclk_2 (pll_0_outclk2_clk), // outclk2.clk
		.locked   ()                   // (terminated)
	);

	ps2 ps2 (
		.clk                   (clk_sys_clk),                                   //               clock.clk
		.io_address            (mm_interconnect_0_ps2_io_address),              //                  io.address
		.io_read               (mm_interconnect_0_ps2_io_read),                 //                    .read
		.io_readdata           (mm_interconnect_0_ps2_io_readdata),             //                    .readdata
		.io_write              (mm_interconnect_0_ps2_io_write),                //                    .write
		.io_writedata          (mm_interconnect_0_ps2_io_writedata),            //                    .writedata
		.sysctl_address        (mm_interconnect_0_ps2_sysctl_address),          //              sysctl.address
		.sysctl_read           (mm_interconnect_0_ps2_sysctl_read),             //                    .read
		.sysctl_readdata       (mm_interconnect_0_ps2_sysctl_readdata),         //                    .readdata
		.sysctl_write          (mm_interconnect_0_ps2_sysctl_write),            //                    .write
		.sysctl_writedata      (mm_interconnect_0_ps2_sysctl_writedata),        //                    .writedata
		.rst_n                 (~reset_sys_reset_out_reset),                    //          reset_sink.reset_n
		.irq_mouse             (irq_mapper_receiver8_irq),                      //           irq_mouse.irq
		.ps2_kbclk             (ps2_kbclk_in),                                  //          export_ps2.kbclk_in
		.ps2_kbdat             (ps2_kbdat_in),                                  //                    .kbdat_in
		.ps2_kbclk_out         (ps2_kbclk_out),                                 //                    .kbclk_out
		.ps2_kbdat_out         (ps2_kbdat_out),                                 //                    .kbdat_out
		.ps2_mouseclk          (ps2_mouseclk_in),                               //                    .mouseclk_in
		.ps2_mousedat          (ps2_mousedat_in),                               //                    .mousedat_in
		.ps2_mouseclk_out      (ps2_mouseclk_out),                              //                    .mouseclk_out
		.ps2_mousedat_out      (ps2_mousedat_out),                              //                    .mousedat_out
		.irq_keyb              (irq_mapper_receiver7_irq),                      //            irq_keyb.irq
		.speaker_61h_read      (ps2_conduit_speaker_61h_speaker_61h_read),      // conduit_speaker_61h.speaker_61h_read
		.speaker_61h_readdata  (pit_conduit_speaker_61h_speaker_61h_readdata),  //                    .speaker_61h_readdata
		.speaker_61h_write     (ps2_conduit_speaker_61h_speaker_61h_write),     //                    .speaker_61h_write
		.speaker_61h_writedata (ps2_conduit_speaker_61h_speaker_61h_writedata), //                    .speaker_61h_writedata
		.output_a20_enable     (ps2_misc_a20_enable),                           // export_ps2_out_port.a20_enable
		.output_reset_n        (ps2_misc_reset_n),                              //                    .reset_n
		.a20_enable            (ps2_conduit_a20_a20_enable)                     //         conduit_a20.a20_enable
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_sys (
		.reset_in0      (qsys_reset_reset),          // reset_in0.reset
		.clk            (clk_sys_clk),               //       clk.clk
		.reset_out      (reset_sys_reset_out_reset), // reset_out.reset
		.reset_req      (),                          // (terminated)
		.reset_req_in0  (1'b0),                      // (terminated)
		.reset_in1      (1'b0),                      // (terminated)
		.reset_req_in1  (1'b0),                      // (terminated)
		.reset_in2      (1'b0),                      // (terminated)
		.reset_req_in2  (1'b0),                      // (terminated)
		.reset_in3      (1'b0),                      // (terminated)
		.reset_req_in3  (1'b0),                      // (terminated)
		.reset_in4      (1'b0),                      // (terminated)
		.reset_req_in4  (1'b0),                      // (terminated)
		.reset_in5      (1'b0),                      // (terminated)
		.reset_req_in5  (1'b0),                      // (terminated)
		.reset_in6      (1'b0),                      // (terminated)
		.reset_req_in6  (1'b0),                      // (terminated)
		.reset_in7      (1'b0),                      // (terminated)
		.reset_req_in7  (1'b0),                      // (terminated)
		.reset_in8      (1'b0),                      // (terminated)
		.reset_req_in8  (1'b0),                      // (terminated)
		.reset_in9      (1'b0),                      // (terminated)
		.reset_req_in9  (1'b0),                      // (terminated)
		.reset_in10     (1'b0),                      // (terminated)
		.reset_req_in10 (1'b0),                      // (terminated)
		.reset_in11     (1'b0),                      // (terminated)
		.reset_req_in11 (1'b0),                      // (terminated)
		.reset_in12     (1'b0),                      // (terminated)
		.reset_req_in12 (1'b0),                      // (terminated)
		.reset_in13     (1'b0),                      // (terminated)
		.reset_req_in13 (1'b0),                      // (terminated)
		.reset_in14     (1'b0),                      // (terminated)
		.reset_req_in14 (1'b0),                      // (terminated)
		.reset_in15     (1'b0),                      // (terminated)
		.reset_req_in15 (1'b0)                       // (terminated)
	);

	rtc rtc (
		.clk            (clk_sys_clk),                          //         clock.clk
		.io_address     (mm_interconnect_0_rtc_io_address),     //            io.address
		.io_read        (mm_interconnect_0_rtc_io_read),        //              .read
		.io_readdata    (mm_interconnect_0_rtc_io_readdata),    //              .readdata
		.io_write       (mm_interconnect_0_rtc_io_write),       //              .write
		.io_writedata   (mm_interconnect_0_rtc_io_writedata),   //              .writedata
		.mgmt_address   (mm_interconnect_1_rtc_mgmt_address),   //          mgmt.address
		.mgmt_write     (mm_interconnect_1_rtc_mgmt_write),     //              .write
		.mgmt_writedata (mm_interconnect_1_rtc_mgmt_writedata), //              .writedata
		.rst_n          (~reset_sys_reset_out_reset),           //    reset_sink.reset_n
		.irq            (irq_mapper_receiver1_irq)              // interrupt_rtc.irq
	);

	sound sound (
		.clk                        (clk_sys_clk),                                               //                    clock.clk
		.io_address                 (mm_interconnect_0_sound_io_address),                        //                       io.address
		.io_read                    (mm_interconnect_0_sound_io_read),                           //                         .read
		.io_readdata                (mm_interconnect_0_sound_io_readdata),                       //                         .readdata
		.io_write                   (mm_interconnect_0_sound_io_write),                          //                         .write
		.io_writedata               (mm_interconnect_0_sound_io_writedata),                      //                         .writedata
		.fm_address                 (mm_interconnect_0_sound_fm_address),                        //                       fm.address
		.fm_read                    (mm_interconnect_0_sound_fm_read),                           //                         .read
		.fm_readdata                (mm_interconnect_0_sound_fm_readdata),                       //                         .readdata
		.fm_write                   (mm_interconnect_0_sound_fm_write),                          //                         .write
		.fm_writedata               (mm_interconnect_0_sound_fm_writedata),                      //                         .writedata
		.mgmt_address               (mm_interconnect_1_sound_mgmt_address),                      //                     mgmt.address
		.mgmt_write                 (mm_interconnect_1_sound_mgmt_write),                        //                         .write
		.mgmt_writedata             (mm_interconnect_1_sound_mgmt_writedata),                    //                         .writedata
		.rst_n                      (~reset_sys_reset_out_reset),                                //               reset_sink.reset_n
		.irq                        (irq_mapper_receiver2_irq),                                  //         interrupt_sender.irq
		.dma_soundblaster_req       (sound_conduit_dma_soundblaster_dma_soundblaster_req),       // conduit_dma_soundblaster.dma_soundblaster_req
		.dma_soundblaster_ack       (pc_dma_conduit_dma_soundblaster_dma_soundblaster_ack),      //                         .dma_soundblaster_ack
		.dma_soundblaster_terminal  (pc_dma_conduit_dma_soundblaster_dma_soundblaster_terminal), //                         .dma_soundblaster_terminal
		.dma_soundblaster_readdata  (pc_dma_conduit_dma_soundblaster_dma_soundblaster_readdata), //                         .dma_soundblaster_readdata
		.dma_soundblaster_writedata (sound_conduit_dma_soundblaster_dma_soundblaster_writedata), //                         .dma_soundblaster_writedata
		.sample_l                   (sound_sample_l),                                            //            conduit_sound.sample_l
		.sample_r                   (sound_sample_r),                                            //                         .sample_r
		.fm_mode                    (sound_fm_mode),                                             //                         .fm_mode
		.mpu_midi_in                (sound_mpu_midi_in),                                         //                         .mpu_midi_in
		.mpu_midi_out               (sound_mpu_midi_out),                                        //                         .mpu_midi_out
		.clk_opl                    (clk_clk),                                                   //                clock_opl.clk
		.mpu_address                (mm_interconnect_0_sound_mpu_address),                       //                      mpu.address
		.mpu_read                   (mm_interconnect_0_sound_mpu_read),                          //                         .read
		.mpu_readdata               (mm_interconnect_0_sound_mpu_readdata),                      //                         .readdata
		.mpu_write                  (mm_interconnect_0_sound_mpu_write),                         //                         .write
		.mpu_writedata              (mm_interconnect_0_sound_mpu_writedata)                      //                         .writedata
	);

	altera_16550_uart #(
		.FAMILY         ("Cyclone V"),
		.MEM_BLOCK_TYPE ("M10K"),
		.FIFO_MODE      (1),
		.FIFO_DEPTH     (32),
		.FIFO_WATERMARK (0),
		.FIFO_HWFC      (0),
		.FIFO_SWFC      (0),
		.DMA_EXTRA      (0)
	) uart (
		.addr            (width_trans_out_address),             //  avalon_slave.address
		.write           (width_trans_out_write),               //              .write
		.writedata       (width_trans_out_writedata),           //              .writedata
		.read            (width_trans_out_read),                //              .read
		.readdata        (width_trans_out_readdata),            //              .readdata
		.clk             (pll_0_outclk2_clk),                   //         clock.clk
		.rst_n           (~rst_controller_001_reset_out_reset), //    reset_sink.reset_n
		.intr            (irq_synchronizer_receiver_irq),       //    irq_sender.irq
		.sin             (uart_s_sin),                          // RS_232_Serial.sin
		.sout            (uart_s_sout),                         //              .sout
		.sout_oe         (uart_s_sout_oe),                      //              .sout_oe
		.cts_n           (uart_h_cts_n),                        //  RS_232_Modem.cts_n
		.rts_n           (uart_h_rts_n),                        //              .rts_n
		.dsr_n           (uart_h_dsr_n),                        //              .dsr_n
		.dcd_n           (uart_h_dcd_n),                        //              .dcd_n
		.ri_n            (uart_h_ri_n),                         //              .ri_n
		.dtr_n           (uart_h_dtr_n),                        //              .dtr_n
		.out1_n          (uart_h_out1_n),                       //              .out1_n
		.out2_n          (uart_h_out2_n),                       //              .out2_n
		.dma_tx_ack_n    (1'b1),                                //   (terminated)
		.dma_tx_req_n    (),                                    //   (terminated)
		.dma_tx_single_n (),                                    //   (terminated)
		.dma_rx_ack_n    (1'b1),                                //   (terminated)
		.dma_rx_req_n    (),                                    //   (terminated)
		.dma_rx_single_n ()                                     //   (terminated)
	);

	vga vga (
		.clk_sys        (clk_sys_clk),                          //        clock_sys.clk
		.clk_vga        (pll_0_outclk1_clk),                    //        clock_vga.clk
		.io_b_address   (mm_interconnect_0_vga_io_b_address),   //             io_b.address
		.io_b_read      (mm_interconnect_0_vga_io_b_read),      //                 .read
		.io_b_readdata  (mm_interconnect_0_vga_io_b_readdata),  //                 .readdata
		.io_b_write     (mm_interconnect_0_vga_io_b_write),     //                 .write
		.io_b_writedata (mm_interconnect_0_vga_io_b_writedata), //                 .writedata
		.io_c_address   (mm_interconnect_0_vga_io_c_address),   //             io_c.address
		.io_c_read      (mm_interconnect_0_vga_io_c_read),      //                 .read
		.io_c_readdata  (mm_interconnect_0_vga_io_c_readdata),  //                 .readdata
		.io_c_write     (mm_interconnect_0_vga_io_c_write),     //                 .write
		.io_c_writedata (mm_interconnect_0_vga_io_c_writedata), //                 .writedata
		.io_d_address   (mm_interconnect_0_vga_io_d_address),   //             io_d.address
		.io_d_read      (mm_interconnect_0_vga_io_d_read),      //                 .read
		.io_d_readdata  (mm_interconnect_0_vga_io_d_readdata),  //                 .readdata
		.io_d_write     (mm_interconnect_0_vga_io_d_write),     //                 .write
		.io_d_writedata (mm_interconnect_0_vga_io_d_writedata), //                 .writedata
		.mem_address    (mm_interconnect_3_vga_mem_address),    //              mem.address
		.mem_read       (mm_interconnect_3_vga_mem_read),       //                 .read
		.mem_readdata   (mm_interconnect_3_vga_mem_readdata),   //                 .readdata
		.mem_write      (mm_interconnect_3_vga_mem_write),      //                 .write
		.mem_writedata  (mm_interconnect_3_vga_mem_writedata),  //                 .writedata
		.rst_n          (~reset_sys_reset_out_reset),           //       reset_sink.reset_n
		.vga_clock      (vga_clock),                            //       export_vga.clock
		.vga_blank_n    (vga_blank_n),                          //                 .blank_n
		.vga_horiz_sync (vga_hsync),                            //                 .hsync
		.vga_vert_sync  (vga_vsync),                            //                 .vsync
		.vga_r          (vga_r),                                //                 .r
		.vga_g          (vga_g),                                //                 .g
		.vga_b          (vga_b),                                //                 .b
		.irq            (irq_mapper_receiver6_irq)              // interrupt_sender.irq
	);

	width_trans width_trans (
		.clk           (pll_0_outclk2_clk),                          // clock.clk
		.reset         (rst_controller_001_reset_out_reset),         // reset.reset
		.in_address    (mm_interconnect_0_width_trans_in_address),   //    in.address
		.in_read       (mm_interconnect_0_width_trans_in_read),      //      .read
		.in_readdata   (mm_interconnect_0_width_trans_in_readdata),  //      .readdata
		.in_write      (mm_interconnect_0_width_trans_in_write),     //      .write
		.in_writedata  (mm_interconnect_0_width_trans_in_writedata), //      .writedata
		.out_address   (width_trans_out_address),                    //   out.address
		.out_read      (width_trans_out_read),                       //      .read
		.out_readdata  (width_trans_out_readdata),                   //      .readdata
		.out_write     (width_trans_out_write),                      //      .write
		.out_writedata (width_trans_out_writedata)                   //      .writedata
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.pll_0_outclk0_clk                             (clk_sys_clk),                                 //                           pll_0_outclk0.clk
		.pll_0_outclk2_clk                             (pll_0_outclk2_clk),                           //                           pll_0_outclk2.clk
		.ao486_reset_sink_reset_bridge_in_reset_reset  (rst_controller_reset_out_reset),              //  ao486_reset_sink_reset_bridge_in_reset.reset
		.sound_reset_sink_reset_bridge_in_reset_reset  (reset_sys_reset_out_reset),                   //  sound_reset_sink_reset_bridge_in_reset.reset
		.width_trans_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),          // width_trans_reset_reset_bridge_in_reset.reset
		.ao486_avalon_io_address                       (ao486_avalon_io_address),                     //                         ao486_avalon_io.address
		.ao486_avalon_io_waitrequest                   (ao486_avalon_io_waitrequest),                 //                                        .waitrequest
		.ao486_avalon_io_byteenable                    (ao486_avalon_io_byteenable),                  //                                        .byteenable
		.ao486_avalon_io_read                          (ao486_avalon_io_read),                        //                                        .read
		.ao486_avalon_io_readdata                      (ao486_avalon_io_readdata),                    //                                        .readdata
		.ao486_avalon_io_readdatavalid                 (ao486_avalon_io_readdatavalid),               //                                        .readdatavalid
		.ao486_avalon_io_write                         (ao486_avalon_io_write),                       //                                        .write
		.ao486_avalon_io_writedata                     (ao486_avalon_io_writedata),                   //                                        .writedata
		.floppy0_io_address                            (mm_interconnect_0_floppy0_io_address),        //                              floppy0_io.address
		.floppy0_io_write                              (mm_interconnect_0_floppy0_io_write),          //                                        .write
		.floppy0_io_read                               (mm_interconnect_0_floppy0_io_read),           //                                        .read
		.floppy0_io_readdata                           (mm_interconnect_0_floppy0_io_readdata),       //                                        .readdata
		.floppy0_io_writedata                          (mm_interconnect_0_floppy0_io_writedata),      //                                        .writedata
		.hdd0_io_address                               (mm_interconnect_0_hdd0_io_address),           //                                 hdd0_io.address
		.hdd0_io_write                                 (mm_interconnect_0_hdd0_io_write),             //                                        .write
		.hdd0_io_read                                  (mm_interconnect_0_hdd0_io_read),              //                                        .read
		.hdd0_io_readdata                              (mm_interconnect_0_hdd0_io_readdata),          //                                        .readdata
		.hdd0_io_writedata                             (mm_interconnect_0_hdd0_io_writedata),         //                                        .writedata
		.hdd0_io_byteenable                            (mm_interconnect_0_hdd0_io_byteenable),        //                                        .byteenable
		.hdd1_io_address                               (mm_interconnect_0_hdd1_io_address),           //                                 hdd1_io.address
		.hdd1_io_write                                 (mm_interconnect_0_hdd1_io_write),             //                                        .write
		.hdd1_io_read                                  (mm_interconnect_0_hdd1_io_read),              //                                        .read
		.hdd1_io_readdata                              (mm_interconnect_0_hdd1_io_readdata),          //                                        .readdata
		.hdd1_io_writedata                             (mm_interconnect_0_hdd1_io_writedata),         //                                        .writedata
		.hdd1_io_byteenable                            (mm_interconnect_0_hdd1_io_byteenable),        //                                        .byteenable
		.hddext_0x370_io_address                       (mm_interconnect_0_hddext_0x370_io_address),   //                         hddext_0x370_io.address
		.hddext_0x370_io_write                         (mm_interconnect_0_hddext_0x370_io_write),     //                                        .write
		.hddext_0x370_io_read                          (mm_interconnect_0_hddext_0x370_io_read),      //                                        .read
		.hddext_0x370_io_readdata                      (mm_interconnect_0_hddext_0x370_io_readdata),  //                                        .readdata
		.hddext_0x370_io_writedata                     (mm_interconnect_0_hddext_0x370_io_writedata), //                                        .writedata
		.pc_dma_master_address                         (mm_interconnect_0_pc_dma_master_address),     //                           pc_dma_master.address
		.pc_dma_master_write                           (mm_interconnect_0_pc_dma_master_write),       //                                        .write
		.pc_dma_master_read                            (mm_interconnect_0_pc_dma_master_read),        //                                        .read
		.pc_dma_master_readdata                        (mm_interconnect_0_pc_dma_master_readdata),    //                                        .readdata
		.pc_dma_master_writedata                       (mm_interconnect_0_pc_dma_master_writedata),   //                                        .writedata
		.pc_dma_page_address                           (mm_interconnect_0_pc_dma_page_address),       //                             pc_dma_page.address
		.pc_dma_page_write                             (mm_interconnect_0_pc_dma_page_write),         //                                        .write
		.pc_dma_page_read                              (mm_interconnect_0_pc_dma_page_read),          //                                        .read
		.pc_dma_page_readdata                          (mm_interconnect_0_pc_dma_page_readdata),      //                                        .readdata
		.pc_dma_page_writedata                         (mm_interconnect_0_pc_dma_page_writedata),     //                                        .writedata
		.pc_dma_slave_address                          (mm_interconnect_0_pc_dma_slave_address),      //                            pc_dma_slave.address
		.pc_dma_slave_write                            (mm_interconnect_0_pc_dma_slave_write),        //                                        .write
		.pc_dma_slave_read                             (mm_interconnect_0_pc_dma_slave_read),         //                                        .read
		.pc_dma_slave_readdata                         (mm_interconnect_0_pc_dma_slave_readdata),     //                                        .readdata
		.pc_dma_slave_writedata                        (mm_interconnect_0_pc_dma_slave_writedata),    //                                        .writedata
		.pic_master_address                            (mm_interconnect_0_pic_master_address),        //                              pic_master.address
		.pic_master_write                              (mm_interconnect_0_pic_master_write),          //                                        .write
		.pic_master_read                               (mm_interconnect_0_pic_master_read),           //                                        .read
		.pic_master_readdata                           (mm_interconnect_0_pic_master_readdata),       //                                        .readdata
		.pic_master_writedata                          (mm_interconnect_0_pic_master_writedata),      //                                        .writedata
		.pic_slave_address                             (mm_interconnect_0_pic_slave_address),         //                               pic_slave.address
		.pic_slave_write                               (mm_interconnect_0_pic_slave_write),           //                                        .write
		.pic_slave_read                                (mm_interconnect_0_pic_slave_read),            //                                        .read
		.pic_slave_readdata                            (mm_interconnect_0_pic_slave_readdata),        //                                        .readdata
		.pic_slave_writedata                           (mm_interconnect_0_pic_slave_writedata),       //                                        .writedata
		.pit_io_address                                (mm_interconnect_0_pit_io_address),            //                                  pit_io.address
		.pit_io_write                                  (mm_interconnect_0_pit_io_write),              //                                        .write
		.pit_io_read                                   (mm_interconnect_0_pit_io_read),               //                                        .read
		.pit_io_readdata                               (mm_interconnect_0_pit_io_readdata),           //                                        .readdata
		.pit_io_writedata                              (mm_interconnect_0_pit_io_writedata),          //                                        .writedata
		.ps2_io_address                                (mm_interconnect_0_ps2_io_address),            //                                  ps2_io.address
		.ps2_io_write                                  (mm_interconnect_0_ps2_io_write),              //                                        .write
		.ps2_io_read                                   (mm_interconnect_0_ps2_io_read),               //                                        .read
		.ps2_io_readdata                               (mm_interconnect_0_ps2_io_readdata),           //                                        .readdata
		.ps2_io_writedata                              (mm_interconnect_0_ps2_io_writedata),          //                                        .writedata
		.ps2_sysctl_address                            (mm_interconnect_0_ps2_sysctl_address),        //                              ps2_sysctl.address
		.ps2_sysctl_write                              (mm_interconnect_0_ps2_sysctl_write),          //                                        .write
		.ps2_sysctl_read                               (mm_interconnect_0_ps2_sysctl_read),           //                                        .read
		.ps2_sysctl_readdata                           (mm_interconnect_0_ps2_sysctl_readdata),       //                                        .readdata
		.ps2_sysctl_writedata                          (mm_interconnect_0_ps2_sysctl_writedata),      //                                        .writedata
		.rtc_io_address                                (mm_interconnect_0_rtc_io_address),            //                                  rtc_io.address
		.rtc_io_write                                  (mm_interconnect_0_rtc_io_write),              //                                        .write
		.rtc_io_read                                   (mm_interconnect_0_rtc_io_read),               //                                        .read
		.rtc_io_readdata                               (mm_interconnect_0_rtc_io_readdata),           //                                        .readdata
		.rtc_io_writedata                              (mm_interconnect_0_rtc_io_writedata),          //                                        .writedata
		.sound_fm_address                              (mm_interconnect_0_sound_fm_address),          //                                sound_fm.address
		.sound_fm_write                                (mm_interconnect_0_sound_fm_write),            //                                        .write
		.sound_fm_read                                 (mm_interconnect_0_sound_fm_read),             //                                        .read
		.sound_fm_readdata                             (mm_interconnect_0_sound_fm_readdata),         //                                        .readdata
		.sound_fm_writedata                            (mm_interconnect_0_sound_fm_writedata),        //                                        .writedata
		.sound_io_address                              (mm_interconnect_0_sound_io_address),          //                                sound_io.address
		.sound_io_write                                (mm_interconnect_0_sound_io_write),            //                                        .write
		.sound_io_read                                 (mm_interconnect_0_sound_io_read),             //                                        .read
		.sound_io_readdata                             (mm_interconnect_0_sound_io_readdata),         //                                        .readdata
		.sound_io_writedata                            (mm_interconnect_0_sound_io_writedata),        //                                        .writedata
		.sound_mpu_address                             (mm_interconnect_0_sound_mpu_address),         //                               sound_mpu.address
		.sound_mpu_write                               (mm_interconnect_0_sound_mpu_write),           //                                        .write
		.sound_mpu_read                                (mm_interconnect_0_sound_mpu_read),            //                                        .read
		.sound_mpu_readdata                            (mm_interconnect_0_sound_mpu_readdata),        //                                        .readdata
		.sound_mpu_writedata                           (mm_interconnect_0_sound_mpu_writedata),       //                                        .writedata
		.vga_io_b_address                              (mm_interconnect_0_vga_io_b_address),          //                                vga_io_b.address
		.vga_io_b_write                                (mm_interconnect_0_vga_io_b_write),            //                                        .write
		.vga_io_b_read                                 (mm_interconnect_0_vga_io_b_read),             //                                        .read
		.vga_io_b_readdata                             (mm_interconnect_0_vga_io_b_readdata),         //                                        .readdata
		.vga_io_b_writedata                            (mm_interconnect_0_vga_io_b_writedata),        //                                        .writedata
		.vga_io_c_address                              (mm_interconnect_0_vga_io_c_address),          //                                vga_io_c.address
		.vga_io_c_write                                (mm_interconnect_0_vga_io_c_write),            //                                        .write
		.vga_io_c_read                                 (mm_interconnect_0_vga_io_c_read),             //                                        .read
		.vga_io_c_readdata                             (mm_interconnect_0_vga_io_c_readdata),         //                                        .readdata
		.vga_io_c_writedata                            (mm_interconnect_0_vga_io_c_writedata),        //                                        .writedata
		.vga_io_d_address                              (mm_interconnect_0_vga_io_d_address),          //                                vga_io_d.address
		.vga_io_d_write                                (mm_interconnect_0_vga_io_d_write),            //                                        .write
		.vga_io_d_read                                 (mm_interconnect_0_vga_io_d_read),             //                                        .read
		.vga_io_d_readdata                             (mm_interconnect_0_vga_io_d_readdata),         //                                        .readdata
		.vga_io_d_writedata                            (mm_interconnect_0_vga_io_d_writedata),        //                                        .writedata
		.width_trans_in_address                        (mm_interconnect_0_width_trans_in_address),    //                          width_trans_in.address
		.width_trans_in_write                          (mm_interconnect_0_width_trans_in_write),      //                                        .write
		.width_trans_in_read                           (mm_interconnect_0_width_trans_in_read),       //                                        .read
		.width_trans_in_readdata                       (mm_interconnect_0_width_trans_in_readdata),   //                                        .readdata
		.width_trans_in_writedata                      (mm_interconnect_0_width_trans_in_writedata)   //                                        .writedata
	);

	system_mm_interconnect_1 mm_interconnect_1 (
		.pll_0_outclk0_clk                                  (clk_sys_clk),                                                          //                            pll_0_outclk0.clk
		.floppy0_reset_sink_reset_bridge_in_reset_reset     (reset_sys_reset_out_reset),                                            // floppy0_reset_sink_reset_bridge_in_reset.reset
		.floppy0_avalon_master_address                      (floppy0_avalon_master_address),                                        //                    floppy0_avalon_master.address
		.floppy0_avalon_master_waitrequest                  (floppy0_avalon_master_waitrequest),                                    //                                         .waitrequest
		.floppy0_avalon_master_read                         (floppy0_avalon_master_read),                                           //                                         .read
		.floppy0_avalon_master_readdata                     (floppy0_avalon_master_readdata),                                       //                                         .readdata
		.floppy0_avalon_master_readdatavalid                (floppy0_avalon_master_readdatavalid),                                  //                                         .readdatavalid
		.floppy0_avalon_master_write                        (floppy0_avalon_master_write),                                          //                                         .write
		.floppy0_avalon_master_writedata                    (floppy0_avalon_master_writedata),                                      //                                         .writedata
		.hdd0_avalon_master_address                         (hdd0_avalon_master_address),                                           //                       hdd0_avalon_master.address
		.hdd0_avalon_master_waitrequest                     (hdd0_avalon_master_waitrequest),                                       //                                         .waitrequest
		.hdd0_avalon_master_read                            (hdd0_avalon_master_read),                                              //                                         .read
		.hdd0_avalon_master_readdata                        (hdd0_avalon_master_readdata),                                          //                                         .readdata
		.hdd0_avalon_master_readdatavalid                   (hdd0_avalon_master_readdatavalid),                                     //                                         .readdatavalid
		.hdd0_avalon_master_write                           (hdd0_avalon_master_write),                                             //                                         .write
		.hdd0_avalon_master_writedata                       (hdd0_avalon_master_writedata),                                         //                                         .writedata
		.hdd1_avalon_master_address                         (hdd1_avalon_master_address),                                           //                       hdd1_avalon_master.address
		.hdd1_avalon_master_waitrequest                     (hdd1_avalon_master_waitrequest),                                       //                                         .waitrequest
		.hdd1_avalon_master_read                            (hdd1_avalon_master_read),                                              //                                         .read
		.hdd1_avalon_master_readdata                        (hdd1_avalon_master_readdata),                                          //                                         .readdata
		.hdd1_avalon_master_readdatavalid                   (hdd1_avalon_master_readdatavalid),                                     //                                         .readdatavalid
		.hdd1_avalon_master_write                           (hdd1_avalon_master_write),                                             //                                         .write
		.hdd1_avalon_master_writedata                       (hdd1_avalon_master_writedata),                                         //                                         .writedata
		.mm_bridge_m0_address                               (mm_bridge_m0_address),                                                 //                             mm_bridge_m0.address
		.mm_bridge_m0_waitrequest                           (mm_bridge_m0_waitrequest),                                             //                                         .waitrequest
		.mm_bridge_m0_burstcount                            (mm_bridge_m0_burstcount),                                              //                                         .burstcount
		.mm_bridge_m0_byteenable                            (mm_bridge_m0_byteenable),                                              //                                         .byteenable
		.mm_bridge_m0_read                                  (mm_bridge_m0_read),                                                    //                                         .read
		.mm_bridge_m0_readdata                              (mm_bridge_m0_readdata),                                                //                                         .readdata
		.mm_bridge_m0_readdatavalid                         (mm_bridge_m0_readdatavalid),                                           //                                         .readdatavalid
		.mm_bridge_m0_write                                 (mm_bridge_m0_write),                                                   //                                         .write
		.mm_bridge_m0_writedata                             (mm_bridge_m0_writedata),                                               //                                         .writedata
		.mm_bridge_m0_debugaccess                           (mm_bridge_m0_debugaccess),                                             //                                         .debugaccess
		.pc_bus_avalon_sdram_master_address                 (pc_bus_avalon_sdram_master_address),                                   //               pc_bus_avalon_sdram_master.address
		.pc_bus_avalon_sdram_master_waitrequest             (pc_bus_avalon_sdram_master_waitrequest),                               //                                         .waitrequest
		.pc_bus_avalon_sdram_master_burstcount              (pc_bus_avalon_sdram_master_burstcount),                                //                                         .burstcount
		.pc_bus_avalon_sdram_master_byteenable              (pc_bus_avalon_sdram_master_byteenable),                                //                                         .byteenable
		.pc_bus_avalon_sdram_master_read                    (pc_bus_avalon_sdram_master_read),                                      //                                         .read
		.pc_bus_avalon_sdram_master_readdata                (pc_bus_avalon_sdram_master_readdata),                                  //                                         .readdata
		.pc_bus_avalon_sdram_master_readdatavalid           (pc_bus_avalon_sdram_master_readdatavalid),                             //                                         .readdatavalid
		.pc_bus_avalon_sdram_master_write                   (pc_bus_avalon_sdram_master_write),                                     //                                         .write
		.pc_bus_avalon_sdram_master_writedata               (pc_bus_avalon_sdram_master_writedata),                                 //                                         .writedata
		.pc_dma_avalon_master_address                       (pc_dma_avalon_master_address),                                         //                     pc_dma_avalon_master.address
		.pc_dma_avalon_master_waitrequest                   (pc_dma_avalon_master_waitrequest),                                     //                                         .waitrequest
		.pc_dma_avalon_master_read                          (pc_dma_avalon_master_read),                                            //                                         .read
		.pc_dma_avalon_master_readdata                      (pc_dma_avalon_master_readdata),                                        //                                         .readdata
		.pc_dma_avalon_master_readdatavalid                 (pc_dma_avalon_master_readdatavalid),                                   //                                         .readdatavalid
		.pc_dma_avalon_master_write                         (pc_dma_avalon_master_write),                                           //                                         .write
		.pc_dma_avalon_master_writedata                     (pc_dma_avalon_master_writedata),                                       //                                         .writedata
		.address_span_extender_windowed_slave_address       (mm_interconnect_1_address_span_extender_windowed_slave_address),       //     address_span_extender_windowed_slave.address
		.address_span_extender_windowed_slave_write         (mm_interconnect_1_address_span_extender_windowed_slave_write),         //                                         .write
		.address_span_extender_windowed_slave_read          (mm_interconnect_1_address_span_extender_windowed_slave_read),          //                                         .read
		.address_span_extender_windowed_slave_readdata      (mm_interconnect_1_address_span_extender_windowed_slave_readdata),      //                                         .readdata
		.address_span_extender_windowed_slave_writedata     (mm_interconnect_1_address_span_extender_windowed_slave_writedata),     //                                         .writedata
		.address_span_extender_windowed_slave_burstcount    (mm_interconnect_1_address_span_extender_windowed_slave_burstcount),    //                                         .burstcount
		.address_span_extender_windowed_slave_byteenable    (mm_interconnect_1_address_span_extender_windowed_slave_byteenable),    //                                         .byteenable
		.address_span_extender_windowed_slave_readdatavalid (mm_interconnect_1_address_span_extender_windowed_slave_readdatavalid), //                                         .readdatavalid
		.address_span_extender_windowed_slave_waitrequest   (mm_interconnect_1_address_span_extender_windowed_slave_waitrequest),   //                                         .waitrequest
		.driver_sd_avalon_slave_0_address                   (mm_interconnect_1_driver_sd_avalon_slave_0_address),                   //                 driver_sd_avalon_slave_0.address
		.driver_sd_avalon_slave_0_write                     (mm_interconnect_1_driver_sd_avalon_slave_0_write),                     //                                         .write
		.driver_sd_avalon_slave_0_read                      (mm_interconnect_1_driver_sd_avalon_slave_0_read),                      //                                         .read
		.driver_sd_avalon_slave_0_readdata                  (mm_interconnect_1_driver_sd_avalon_slave_0_readdata),                  //                                         .readdata
		.driver_sd_avalon_slave_0_writedata                 (mm_interconnect_1_driver_sd_avalon_slave_0_writedata),                 //                                         .writedata
		.floppy0_mgmt_address                               (mm_interconnect_1_floppy0_mgmt_address),                               //                             floppy0_mgmt.address
		.floppy0_mgmt_write                                 (mm_interconnect_1_floppy0_mgmt_write),                                 //                                         .write
		.floppy0_mgmt_writedata                             (mm_interconnect_1_floppy0_mgmt_writedata),                             //                                         .writedata
		.floppy0_sd_slave_address                           (mm_interconnect_1_floppy0_sd_slave_address),                           //                         floppy0_sd_slave.address
		.floppy0_sd_slave_write                             (mm_interconnect_1_floppy0_sd_slave_write),                             //                                         .write
		.floppy0_sd_slave_read                              (mm_interconnect_1_floppy0_sd_slave_read),                              //                                         .read
		.floppy0_sd_slave_readdata                          (mm_interconnect_1_floppy0_sd_slave_readdata),                          //                                         .readdata
		.floppy0_sd_slave_writedata                         (mm_interconnect_1_floppy0_sd_slave_writedata),                         //                                         .writedata
		.hdd0_mgmt_address                                  (mm_interconnect_1_hdd0_mgmt_address),                                  //                                hdd0_mgmt.address
		.hdd0_mgmt_write                                    (mm_interconnect_1_hdd0_mgmt_write),                                    //                                         .write
		.hdd0_mgmt_writedata                                (mm_interconnect_1_hdd0_mgmt_writedata),                                //                                         .writedata
		.hdd0_sd_slave_address                              (mm_interconnect_1_hdd0_sd_slave_address),                              //                            hdd0_sd_slave.address
		.hdd0_sd_slave_write                                (mm_interconnect_1_hdd0_sd_slave_write),                                //                                         .write
		.hdd0_sd_slave_read                                 (mm_interconnect_1_hdd0_sd_slave_read),                                 //                                         .read
		.hdd0_sd_slave_readdata                             (mm_interconnect_1_hdd0_sd_slave_readdata),                             //                                         .readdata
		.hdd0_sd_slave_writedata                            (mm_interconnect_1_hdd0_sd_slave_writedata),                            //                                         .writedata
		.hdd1_mgmt_address                                  (mm_interconnect_1_hdd1_mgmt_address),                                  //                                hdd1_mgmt.address
		.hdd1_mgmt_write                                    (mm_interconnect_1_hdd1_mgmt_write),                                    //                                         .write
		.hdd1_mgmt_writedata                                (mm_interconnect_1_hdd1_mgmt_writedata),                                //                                         .writedata
		.hdd1_sd_slave_address                              (mm_interconnect_1_hdd1_sd_slave_address),                              //                            hdd1_sd_slave.address
		.hdd1_sd_slave_write                                (mm_interconnect_1_hdd1_sd_slave_write),                                //                                         .write
		.hdd1_sd_slave_read                                 (mm_interconnect_1_hdd1_sd_slave_read),                                 //                                         .read
		.hdd1_sd_slave_readdata                             (mm_interconnect_1_hdd1_sd_slave_readdata),                             //                                         .readdata
		.hdd1_sd_slave_writedata                            (mm_interconnect_1_hdd1_sd_slave_writedata),                            //                                         .writedata
		.pc_bus_ctrl_address                                (mm_interconnect_1_pc_bus_ctrl_address),                                //                              pc_bus_ctrl.address
		.pc_bus_ctrl_write                                  (mm_interconnect_1_pc_bus_ctrl_write),                                  //                                         .write
		.pc_bus_ctrl_writedata                              (mm_interconnect_1_pc_bus_ctrl_writedata),                              //                                         .writedata
		.pit_mgmt_address                                   (mm_interconnect_1_pit_mgmt_address),                                   //                                 pit_mgmt.address
		.pit_mgmt_write                                     (mm_interconnect_1_pit_mgmt_write),                                     //                                         .write
		.pit_mgmt_writedata                                 (mm_interconnect_1_pit_mgmt_writedata),                                 //                                         .writedata
		.rtc_mgmt_address                                   (mm_interconnect_1_rtc_mgmt_address),                                   //                                 rtc_mgmt.address
		.rtc_mgmt_write                                     (mm_interconnect_1_rtc_mgmt_write),                                     //                                         .write
		.rtc_mgmt_writedata                                 (mm_interconnect_1_rtc_mgmt_writedata),                                 //                                         .writedata
		.sound_mgmt_address                                 (mm_interconnect_1_sound_mgmt_address),                                 //                               sound_mgmt.address
		.sound_mgmt_write                                   (mm_interconnect_1_sound_mgmt_write),                                   //                                         .write
		.sound_mgmt_writedata                               (mm_interconnect_1_sound_mgmt_writedata)                                //                                         .writedata
	);

	system_mm_interconnect_3 mm_interconnect_3 (
		.pll_0_outclk0_clk                             (clk_sys_clk),                            //                           pll_0_outclk0.clk
		.pc_bus_reset_sink_reset_bridge_in_reset_reset (reset_sys_reset_out_reset),              // pc_bus_reset_sink_reset_bridge_in_reset.reset
		.pc_bus_avalon_vga_master_address              (pc_bus_avalon_vga_master_address),       //                pc_bus_avalon_vga_master.address
		.pc_bus_avalon_vga_master_waitrequest          (pc_bus_avalon_vga_master_waitrequest),   //                                        .waitrequest
		.pc_bus_avalon_vga_master_burstcount           (pc_bus_avalon_vga_master_burstcount),    //                                        .burstcount
		.pc_bus_avalon_vga_master_byteenable           (pc_bus_avalon_vga_master_byteenable),    //                                        .byteenable
		.pc_bus_avalon_vga_master_read                 (pc_bus_avalon_vga_master_read),          //                                        .read
		.pc_bus_avalon_vga_master_readdata             (pc_bus_avalon_vga_master_readdata),      //                                        .readdata
		.pc_bus_avalon_vga_master_readdatavalid        (pc_bus_avalon_vga_master_readdatavalid), //                                        .readdatavalid
		.pc_bus_avalon_vga_master_write                (pc_bus_avalon_vga_master_write),         //                                        .write
		.pc_bus_avalon_vga_master_writedata            (pc_bus_avalon_vga_master_writedata),     //                                        .writedata
		.vga_mem_address                               (mm_interconnect_3_vga_mem_address),      //                                 vga_mem.address
		.vga_mem_write                                 (mm_interconnect_3_vga_mem_write),        //                                        .write
		.vga_mem_read                                  (mm_interconnect_3_vga_mem_read),         //                                        .read
		.vga_mem_readdata                              (mm_interconnect_3_vga_mem_readdata),     //                                        .readdata
		.vga_mem_writedata                             (mm_interconnect_3_vga_mem_writedata)     //                                        .writedata
	);

	system_irq_mapper irq_mapper (
		.clk           (clk_sys_clk),                //       clk.clk
		.reset         (reset_sys_reset_out_reset),  // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),   // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),   // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),   // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),   // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),   // receiver5.irq
		.receiver6_irq (irq_mapper_receiver6_irq),   // receiver6.irq
		.receiver7_irq (irq_mapper_receiver7_irq),   // receiver7.irq
		.receiver8_irq (irq_mapper_receiver8_irq),   // receiver8.irq
		.receiver9_irq (irq_mapper_receiver9_irq),   // receiver9.irq
		.sender_irq    (pic_interrupt_receiver_irq)  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (pll_0_outclk2_clk),                  //       receiver_clk.clk
		.sender_clk     (clk_sys_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (reset_sys_reset_out_reset),          //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver9_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (cpu_reset_reset),                // reset_in0.reset
		.clk            (clk_sys_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (reset_sys_reset_out_reset),          // reset_in0.reset
		.clk            (pll_0_outclk2_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
