��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�v���"ӔA����l�����;[�"�9����>�p�[g5~ď8&��v�<d.��"J9qZ\�ѶG�k_������<����5�9o�b�+�%M�VRA� b4?4N�P��A-Y��6�����_
���Jzo�*�^���jR�eU_.䞌km>�ӎpx�2��Ɉ��p�~�/���4�¼�C(�����*���"I�E�ʪ���k��Y�3��;��l���g+��J��"׮o[�~�'��o���I��|�Ĉrޏ�v�����ى,mh�xr�\�����#˙�t�m�,"�%��G�6%���z�Ml���.� G�M�n��*��@��I��}�1+�tw�l����M���a�1}�p����o��'M�։]��`i`�j�o���<��4���j\�ߖ3�;d����z(���O�GV;"<��a�O�c^�(�ӝ��������o)����ۊ��"0aY|����~���K�Ti����
�T_p����>Q.��.9W�v������F�ad��5 �+�����1�,7�<��s?����r+P��äy����E�����Q�cC����#��$z��:i}��De ���T�^�u��?��k<m]�*������ʮAݏ* B�l�dC}��1��#��oK��jK��E�C�5Ö��ee��z~p��[
�ڝG-�O ���9g�=�y��v_�6���>/W�:�{�j�olE�q�G��;�ig]}"O�/$�B����$mW5���ĸ�B��u1N�^c<��F�-��.\�և��(9�4G1�v7���pF����]#a�A��S����.dT���	������<"Y�� �B�OTZ��.�N���=Ȏ�5U 0ۖ�tBlO��k�k�����Q��FS��h:�-����ԳaR�[��g�]�+��D^�@U�]��e�)���O�X&!�&EjL��)*%��K��L�����3��79�l]�8 ��_��	�ޔ��mE�J�e���[�Ҟ?Vԭ�F��	�צSt�n��K8Ē�;�@|�v'3p���N���jw�*;�AF�JL������:i=��r�� �[&򼡳'$�|k��ӟP���Z�J�S�]O�y������'�w`��c�DUU2��-csGꞜ�`y����Bj����s��CTN�s[�:E��7r�Ϻ�w̉�V/���lAh(Q��x�'���ˇ�W����X:1l�Lx)e��Ĩ���id$��rzҲ>��\���R���[��}�.j3�J�����T_���u?���ISsF�Cn �������_��v�)�?>(��y���OجJo��T`}�g�<c�(�M�2�D'�JIȨ1�7�x�l7S��Sř����=��1���+B&�g�7`�)el��II�Ь{��	(X�b`�����ɥE���/���8���vzQpj,�J����O���Q:|Zj�;��.,�#>��?��?�K+�����
�]m=^3PtK��6D��~�%g�4��rS���D��nB<~�I'�H٧;��߇�}���lm#�ԢM<��|A*~��Y�6o�:��&��֚=Z�`�3��5u�E.�QX]�2?��$��Hc-��9,��F��jұ��j�U���F	��� ���M�l^����4�M�������yK^��z�kb�����^����)TE̿���=��%��\���mP���h�<e��2u�wk��:W �&��2���"�1u�v�ӫWYb��@'�N {g���?K) ��Њ�;XL���v�x��-�ɬq�������
 ����"|�fE�9ވWYmw�e���K^KU�=���w���8�=���D�.�%_q�1�2�I"z��j���Q�[�+��}��=�I_��1��=.�ˋ5� WQ�Fe�_b���&
t+ԩ n�������()J'N� L�~|�"�0ՠ���-[�F�1�r)�jS�