��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չk��n�AEfs"�mh���Q��w6Ww��e���mJ�?��ZWjy<���7x���]4���f�m��IȨ�`�43Fy b�G�>����5'-��k����`��|�ү�9������sa�y5-�=��׽u����kh�8=�����=�� �y�z��_�*rR�%�Y�|3'Z`�pjc�g#Q�c��;Sa9@bʑ�|v3	�3�w�p0��E�m�
���S��Kf"X}g?�)ׁ�v4��f �0S�!}�ŤQ@8���֗������]��A�������d�WT���!	����4�9B��T�����߷��1� �/�>�i���jzuM0W	�M�0m:�0"M]�_��t�?�"JC�;��VVv$wVψ���zV��j�_�ؾ��9�+����*�aɸ	��z�p�y��S��I�έ�A���I�
6U^�W�DW(4Q��&��Sa�MȃaJ�I�jf��?��;�b��� ��յv�[]�݂x�� X��`�iG�D��Me�e�Ιf���#�)�v�Z|8�F�]2p�|�{�!r�/��7I�M�<p��}�m&n��!qi艤�v��dC�r���q5�\���<���w���?��f��b�z����:��}@��%ߊ)7|jwa��Qt��b�>+߹���~ŗPR�o3��Wn�����l��7�
��Q�*��9�����|�q:����1�:o�>�c��՝R�.�@&H�~�
G5wO�jZ�;�����:�*`H�O(!_�����_~L��مaH�p��Ǜ�E@0V�R<�vy	�ló��������7{>pCMU���kmu[���,�iˋ(�ι:�!��
ܴ�}�o�����,v{���s�Y�U�/�ʝ��4�aA(��G�鴊�ˑ�-�b�1RayÜ�L�Y�?Z!�TF�%�]WRݳ��z���6.9�&�h�Hc88
=�z�v���&)�2P��@j&(��M>�ϰ�ϩhI�X��U.��ɢe��� �y��q������]_B�X�b�9%��Q��)3X���Z��?�2I�c�f�d)�.�� s�����vS;���M���eN����� z8����x
�� ��B����P�ң��1���E �u�)Mw�+�[��[�:m�y�+-�p��~�KP�s�vB��Ur9bM��˟L1V{��=���z4_����Q}���c�wc���b#�:-r���
�Nv�e(�t�.��k�Vx�q�WI!��1]"��ReK����-�q~$
>�)�]_T�7(i5�^���4"���%Hҫ���T������'���`L/���bn�P"��X�#��C*An/BK��ͺ�8 �h�`i���e\�ʅ��]���e�|4�#.�Z��6��%$\��K����3~�a"1 p�C*����Ի�C]��.NN�ؖrAA���]�b�;Fl�S�X�:����~�zQ���5n�� K�Vk�\�P}Ol�+j);H��iMH��4��;(?��95�b����)?LB;�(,�/y2��͵L�����N�|8�K���HP�K��B���1�YG��.d���+;�)50���p�ʤ-	��yS)� �2�l����D|*�.3�����y��px�(GMI;D4ݧ��)D��[���� ��	j2H9xαL�rc̓/ȃ7E�?ʉ7�:���吶"��Fړ��Vy�(�b=��Ϙ\��PffK�E��o��n��	�N쫹�F+�#b���E�Ԛ�'�I��!ҿ�4"���M��D�<*��͐��� 8�r�BA���f���ڋ���'����sY���$�3����U�04�W���oqҶJS8-o�씀\�	�zu;��ќ�L����<�����T��4����N;۲�v�ݬg3�(��-A���M�\���5��m�'��lxnj0f��c�-_^v�ʶ�V�_+�d��l&}k���ᢱ��Y쏚J�>�)�F��4�#���'��B�[7�>��j��m�@�g��N\�K(j:�q���"i0D���qATi��d7l3n����tu6�3��/u���̼]ya�M$�.��d �n�����{��7�:l|kwL�Rf���G��ڣJ��ub�zWt�6`X�5�-gt�@6Pn�'�n���	T��s�;����v�Fu�C&�H�;�QI��p���KͶ����􎶏����Jp�O��w(|�o��	Dz�� *  [�EhfE�O� �={:]��#��-sA�t��|T9r+d��'���$*,���ho�;4�̓��B\FRE��[��#�^������A"���.wKB�f��x�'�������x&�r��޽�.�? �b��������m���<��ā��7���SN.�����¹eFAf�)O�y���X�$�:_w�m�K9�c�hf����_����KZ�����൅�N�w��D�C<Î������vD���w�\?�M�<��m2�e����k��5P̒�
:��C�o�A�#��i YO����x� G��[�����U!b[�����|�i��b��N�}kmtA<�� �����4`�c���t��J�T��v�R�cY��gͥR]'�5���f��VV?5�!icD��i��e6/���~ál(��]��=�?H��9S��b�à���v �'����F��.-���_m�O��9��Qϝ�ό�+��
�^�Y�d7�x�M}�.-�?�2EQ $��\��!�v���5��UР�4V铼�{`
z'`����[����s��m�1��J9���5[n�73�ܔRq�nN�uW2) ����A�P�Y���=�eDp@&ak�4pUe`H��A�V.������g�7��O?N�^�Ú��$e�O7�!�}H��:2��虴�?@}I�d���=m�!���ؾ�02��_��k��3��t�����&��]�&�H�ۈ�P�O.�����.�_�(hB�0F�g�o?��&�2gb-)��o��lҋB*^�:/a��Fh;t�y����(y�����%o�wp��'vp���f�������c�?�G����+{%+��0�g�����e���ѣ+��s#9F���i��a��͉pq\}$��9Nߦl��e���%bw����Y�w�V�q���{�cz;N#��R��lꪫ�5F��R�]I��  �����E`Hj��T%UJ��ڹGs�պ��k��L?E��X�"�U)+&L8(���ܲ���&�h�,��D���w�ʘ64E��sWOa[ŕ�.Oe`�X�Y�&�k�Y���`�A<a�~ɛȜ�a.����y6W��>ŵU@t�׽9M����4�u]krސ��1U9wg���r���"����"��Z>>4-�ǝ���%�7H���
ߎcl�r�~��������,UԄ�2B�ԭ���Y�ws/�@�᠈Zf��X�� ��1�c�)��TO��)eb{�A ����+U�F�Y�R���jwtY�o�ϥ����<�t��0۳b�*�\�Rp�#���΅r�	<b7L��n���Ϝ��e�B���j�Wx�D-=��%�G>D�ʝ掗u����>�1ڍ*�kL1`��<���0�(L��7Q��4��?	���/u���p��������nqB�,"�`[
�z�zH��P�@Յ(� ��!4��J�`~
v����y�&�t��X�������P����@с�4�ݚ��2�!�sB�m�|>H�R�|O��uW�ad���i��n�r�o���5/���9e����4ė\�_r ��&�TȊ0���*DY6�"������bZV�8���"����L��$4Z+�e�.��WoG �]�m�V9:�T��jOV=Dc/*�0�sR�r/ius��L�SR��/���=fY<�]&ز�tCV\����;%�<#;aO�@���� i9�eWlT�?�C�P��߇`*��T߿a5������jPC�k�F��9��E�Y-���Hz���#g���(%ŏ�ֆۏ	�]�-�t�9����2���Y��c��S���"��F��ѷi�L���D��	�V�Y��R�ۉ��;d2d�-'��)�Sȋ����
D��*o���,�1
*`$^�Ĕ]�Kg�4�t�M�A�dM,v$�7�ȜWN�oV���a\��J�(13+�YW����9���9b�_��3C��|���������h�������yVA��7ü+��S�f�X�.[B*]�L}r�-q)��<�n�Y�݌ڙ/�Ί��d\�@���dӽ��A�]�U#��	qBUј�d��q�����d��͗>#�ğ��17K0��oA��Q����ö���N�#�H�s(�B�S���1�,Gė	b�8�=���^e�f}�: ��o�lr� ��
�4w��V��)�	���͙G�}U F,/j�Y7������{OnEң�F>2L�<\V+
��HR�
�`�M��e��:/�����~Y��D�ݿ������K��͂��x���Y�t�Z�V��#�	���(�0>�	1���>lX�G�*�*�\Q��#�*�O=A�O��3(Ѱˮp�v4���{�w��϶���r�F�]��x���l��Ay�d�q|P�O�]��(j��� w���h��L�	�mZ5ؐÇ����hơ�I��Q���~����$ʁ�WL�a1�i�'�1��Ꮢ%5�ַp�A%+��:5���')�z���x~,{"����������|�^�7�*��T?:^��]w��D5/��bJ.�I����BJ�$�	�b�|�p�4r2� �v��j��H�	[x����N8�JO�O��w<�����Q%l�����ғ4��_���7Q@����o.m
�mc<g�����D��6�*��3g�V�Ŵ�?��	�rX��@ߗ��0���� ��Ϧ����I����?} w���x�Ǿ��-�rn�[��'�p6�o\��O3*�g1��/��Fp�r�Rb��5�z_d�t_��wOoS��j��)��Q�JYj�qvٔ��JMw��]��SLY,��Ċh��mDZ�0�[�Զ��;������B�&��KR�y�g�o�t�lz��E���2a{v�