��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�M��8W�Bek�9|��9��O�:���w����,r�R[��3'?kE�v�b!�H�c��6����0�
��P�p�LηQ�,x�LzK�_��x�S���� F�|"z��Sԧ(Tt%��`���sօR�s)3`���\�z��e�0�c������=V��r�C�b�oH�K��v	�أ��햶1#bV����C��?����ϔ�!2�a���(�Ag�h� (�\�����4яЦ�Vo�]������dX�>�8�%�#R�N�v�~���h�)� �^��d����~����3o��>�Ϯqal��U���8Dy�#M�!��]j�;c×���vo�U�ǌlfDŘ��d�0$璑Kk@x#X=m?��3�V��ՙD�m�i�:{.��;(�x�K��A=&E��:䳕+�0[9����軑���~K%�$�*��k�/�`7G���m1+�_��M��#p�[e̫�+Pd�i�:]7ȳ��|��L�0Y�;�m(JJCN\!��CG��/�0��`Za}��+G�3�by~��-� x�
}�!k@����s���7#9;Ҝ��r�XT�`!�-�ۀu�lw��/u�B��qy����]�`X���N4oގT���UzUe�"d��fJE��HBA���$ <����]9�V�1D���T��=
6��;ε�iw�ߵH��	�t5���pd�"�\sUql��k�<J���uTU�彎_�N��oo��\��>���Q09��}Y{#�[>���X���_��I�f��5l���Rȑ���?�"_W�� ���i�(���_�&��,�P>E�"+ž'M �㡼�D�c@����{	�~���gÔ�$m�NOc46Yx=�m����Y2♴E[���ZZJD�	q�w�|#͠�k��^�s0����#�@j0�k"L�a|2��{�N���/��1J�\:�3�=;�v��w��֞���8>TBA��x)ι��⥬>-���ސ\���-��W`b�xeZ?����yp8�@u��}�n�=tA�ո�����M�B���͢�69��b��r���ک�������V�W��Bl���E2��%) C'nZf醷����7�/Z�y���8��0E}ҡ�UN1�!�͎�ȼn�4�A�h�9O�� �m87�M�Ƅ��,%�>Z�C����0bP�^u�u����6��!H��� ����3B���;��b���~��a��W6�)Iʄ�=�������(�$n���/��'�`aF�B0Bnu��r��e���On�a�L*���&E�,{ݫ�a�v)f���W�՘�enpY� \��/�J���,�kC,��� R�
��j���Q|, ��lE�Tz�Ṃ�y�u�6�)�@�3Eќj�'�n݁n@7QƵ�wd||��}�5��R��}x@�|��r���Ɉ�&9Qd??�e\�_��ȇ��m��=sH�2�-%�������0��.��W����L����'�P\XF�e�=&�r���
�,<��Hh����3'���P�/0��
�5E�9�ۢ�^�c<���Ǽ���P���k��B��Z�L�������ҏN�)	v|���
�ڳ��ҫ�x �wȵ���w�jJ�����i���C����^yv����H�)�rT$�aB��@+�^��*� ��{b5�"*�Jд�%���C�����􈍪�B �;@�k���ij�G^�/�qZ�
�V{L1�<S8ʙ|h>�=�l�w��g}�#x����w�o�����3�c����<��ƭ�b|A[M��묉�����Q^�i�D\�C�&�5(�#�"a2��U]�$��{Sb<bw�$O���Fj���U�3`A�u�uJ�J�9v�>iT^L[-�R�$#����=r�P�&;&>G�\֧��l�X�wO�2�:�.G3ۃ��S���7�����`I[�I�oN-��8��#?kf���B��g�x�j'���>"�i�|m\�F���^�d��2�:���
;�NE���H��a뫏R�s
���ZI)2��Up���5���0Ɂ�P�|�x8g	���2飜�P�W�q;P�q�J�6��sB��jm�48ٙ��je�С�Jǟ���v�B��K y���`u�m��q���ĸ��;�F":u�9ۜ�ֶgZq��H����\Y�p�+��L��)�+�Q���c�����_�v���HO���H�0�׀��3��F���Yv`����
u
^��s�Do�8��dkf&���czVe��(̥"�< K!���H��n�\c�eQi}m-�i֗���:���S:R�K_T�5�s}���[6TX�8�c���t�(����q�M^d�M���x����Z��0v5�K�#b��Æ�`��E��;�j���f�nB�Q�9�-\�R�}�?��b�:�6^�SZ�4�T����=�[�3 В�S(�-��½v�F8�(C`����>�{�C�H�����<(v�/��e\��&̀@�ABFbBi�of��=�o�r��������f�b\mBk�I�,�/�s��ꋾ1�s�HХ� 8q���Z ).�N��h��2,'����:� 5a�<��������Y�'�%��W[eG�Ґ���`2��z�"��.=ȾܬV���PѪ�Ԙ��7��2=����^,�^�]�o�:���	?eLBG��ZM�у>�yG�����2
