--===========================================================================----
--
--  S Y N T H E Z I A B L E    2K Synchronous RAM Module
--
--  www.OpenCores.Org - September 2003
--  This core adheres to the GNU public license  
--
-- File name      : blockram.vhd
--
-- Purpose        : 2KByte Block RAM instance
--
-- Dependencies   : ieee.Std_Logic_1164
--                  ieee.std_logic_unsigned
--                  ieee.std_logic_arith
--                  unisim
--
-- Uses           : RAMB4_S8 from Xilinx Web pack ISE 4.2.03i
--
-- Author         : John E. Kent      
--
--===========================================================================----
--
-- Revision History:
--===========================================================================--
--
-- Version 1.0 
-- John Kent - 6 Sep 2003 - Initial release to Open Cores
--
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library unisim;
	use unisim.all;

entity block_ram is
    Port (
       MEMclk   : in  std_logic;
       MEMcs    : in  std_logic;
		 MEMrw    : in  std_logic;
       MEMaddr  : in  std_logic_vector (10 downto 0);
       MEMrdata : out std_logic_vector (7 downto 0);
       MEMwdata : in  std_logic_vector (7 downto 0)
    );
end block_ram;

architecture rtl of block_ram is

   signal dout0 : std_logic_vector (7 downto 0);
   signal dout1 : std_logic_vector (7 downto 0);
   signal dout2 : std_logic_vector (7 downto 0);
   signal dout3 : std_logic_vector (7 downto 0);

   signal ena0 : std_logic;
   signal ena1 : std_logic;
   signal ena2 : std_logic;
   signal ena3 : std_logic;

	signal we   : std_logic;
   signal reset : std_logic;

   component RAMB4_S8
    generic (
      INIT_00, INIT_01, INIT_02, INIT_03,
	   INIT_04, INIT_05, INIT_06, INIT_07,
	   INIT_08, INIT_09, INIT_0A, INIT_0B,
      INIT_0C, INIT_0D, INIT_0E, INIT_0F : bit_vector (255 downto 0)
    );

    port (
      clk, we, en, rst : in std_logic;
      addr : in std_logic_vector(8 downto 0);
      di : in std_logic_vector(7 downto 0);
      do : out std_logic_vector(7 downto 0)
    );
  end component;

begin

  RAM0 : RAMB4_S8
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map ( clk => MEMclk,
	            en => ena0,
				   we => we,
				   rst => reset,
				   addr(8 downto 0) => MEMaddr(8 downto 0),
               di(7 downto 0)   => MEMwdata,
				   do(7 downto 0)   => dout0(7 downto 0)
	);

  RAM1 : RAMB4_S8
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map ( clk => MEMclk,
	            en => ena1,
				   we => we,
				   rst => reset,
				   addr(8 downto 0) => MEMaddr(8 downto 0),
               di(7 downto 0)   => MEMwdata,
				   do(7 downto 0)   => dout1(7 downto 0)
	);

  RAM2 : RAMB4_S8
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map ( clk => MEMclk,
	            en => ena2,
				   we => we,
				   rst => reset,
				   addr(8 downto 0) => MEMaddr(8 downto 0),
               di(7 downto 0)   => MEMwdata,
				   do(7 downto 0)   => dout2(7 downto 0)
	);

  RAM3 : RAMB4_S8
    generic map ( 
    INIT_00 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_01 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_02 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_03 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_04 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_05 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_06 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_07 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_08 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_09 => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0A => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0B => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0C => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0D => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0E => x"0000000000000000000000000000000000000000000000000000000000000000",
    INIT_0F => x"0000000000000000000000000000000000000000000000000000000000000000"
    )

    port map ( clk => MEMclk,
	            en => ena3,
				   we => we,
				   rst => reset,
				   addr(8 downto 0) => MEMaddr(8 downto 0),
               di(7 downto 0)   => MEMwdata,
				   do(7 downto 0)   => dout3(7 downto 0)
	);

my_ram : process ( MEMaddr, MEMrw, MEMcs, dout0, dout1, dout2, dout3 )
begin
		   case MEMaddr(10 downto 9) is
			when "00" =>
			   ena0  <= '1';
				ena1  <= '0';
				ena2  <= '0';
				ena3  <= '0';
			when "01" =>
			   ena0  <= '0';
				ena1  <= '1';
				ena2  <= '0';
				ena3  <= '0';
			when "10" =>
			   ena0  <= '0';
				ena1  <= '0';
				ena2  <= '1';
				ena3  <= '0';
			when "11" =>
			   ena0  <= '0';
				ena1  <= '0';
				ena2  <= '0';
				ena3  <= '1';
			when others =>
			   ena0  <= '0';
				ena1  <= '0';
				ena2  <= '0';
				ena3  <= '0';
			end case;

		   case MEMaddr(10 downto 9) is
			when "00" =>
            MEMrdata <= dout0;
			when "01" =>
            MEMrdata <= dout1;
			when "10" =>
            MEMrdata <= dout2;
			when "11" =>
            MEMrdata <= dout3;
			when others =>
            MEMrdata <= "00000000";
			end case;

         we <= MEMcs and (not MEMrw);
         reset <= '0';

end process my_ram;

end;

