��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��ՉU��e����_X������pbۣ�"c	�l�P�� �p���cx��PI_T\��Z]M:��M�l��D�LQ�)��p^���E��ӷ�mı���yM��s ��$i�m�<8f��!u���2`6J#y_��>��^J^��`�/.�T���*&��B:�|/�?���BM����um1�k���t��d�=�,o�r�KHW������,��ޝ��.ݷ�����u�P��

��g�Zn�ۗWHݐ��#�A����CJ�M�ԙI؎�"p�����:nn���	W˦2-�vrogV���Ѥ����I�����������Ԙ˧c��0�d�M{��5�:���#ԟ�q���T�R�̚��K}��j@ҹ#������*������}f<,��E�c���{�?��B �	 �ܚ[q&�^����|��
���l<ıY� ��O���d��1'Sv ��`~>o��F����F8�A'��-W��!�� ��U͑/�lAS�f�> �e'ƴ�����%�mR�1�/��q�Bc:��L�ԋ��I�٬U��o26,�ġ�y���+v�4��h�ږ?�*�{N���R���i���`�z��-.RT����J:�g��pŢT)XóL��@0~+�c#g����æ��W�*�z���VA�����3����^���r>b.l�o�?`S�#yȞ8�3����O��Q��!g���W�#��Q�����9�q�m�H��hSLy�����zc޼$p���'Da����n�	MEm�I�#M�^g�-ʎ�m�s�+0�y�D��i���������r�sU��h�G9Bly
5t��f��,�ʑN7��J�ҋAa+l�#~]�g���E hc�t�/\�+�UCJ�����'��	�����,µu���U�5��o��ɔ�tW޺��T٫�Xlke~@8��Wp������5@\)-l��p��pC�Tƛc^�xg��! �n�.�7E����6;�3�)�V�Y��1��.0�)��q�ðH2�@����|�Dxuh���Y�E��	꜂�g�I�b!���,5�)x�(�-��9��n:`A�<K%;����醟�c�d��q��(j9�2�mK.e3V1o\F�O�zQ���$4m��\V�g�T6����oWWu�cC��yXM�\�����_���T���Z��|Y���o�q��@��lCK�z���y ����|e[C��޾�U ��uu�ȉ�Ƴ�`鍩�| �B�V�)��"�"�>�v/�]�;�� ��̲�A�n�L�h5NE�"�b_� յ��)9g�M'o�QfX��0Vm�G�����r�a�� G��	?Qp�si6�p�t��ό�)�� ���l���Âx�8����q�̿;�������z] n�S��Q����ʉ��x��g~��6��p���<�-��'9�AD���W��3
A�㍌H�rur�#K�M@H���kF,:�� Lj���e>p�g��Q�����?�]�-*!��{}��(@����,�L")`�ExD�#��]��kٲ�7�4v�qӣd1	����0�w=
=4��*���5����\ơ��� D��
�\gb�	�n��(�5���q���5��N�J�I��׵/��R����m/Q%ԼjMk����`�l0%n���5P����)�H��c �i1	~O�w3ϫ��8�ٟ�
����>N����"�Ɋ*�k��v�
��{�0�@�h���vKJ�o
�� ��2l~p3a�g��<���7)�%���Aa?���?��uj�u.t�����z�2<���xc-b�&*�������Dvǳ���HKgo��$Me��4B��ly�Gv��D�8�Hdn�)h�j���TLm�)����x,�9hz�`�����l2�OR�2��}��s����QRs��#Q�i��2��h�#&��΀�T�{XjW���	�C�қ��[����;l �	�-Ÿ�`�|J[y!�h�/�v?j��pȞ?�B%,❦�m!K�_�V�R(ǒw�2�i4�,u�'%o��pMn�doZm,?�q3̶���c��5������������TA:=�q�H/.J���t�v�H!��Z�bЋ�� ��0��%D���#� �݇)I�3r����� �[����~��/T-\��~$c�/��x�+�Q�������U��_"���e�Sb:r�<W@�x�B�k!j�J���)�#����A��g��% ƺ��\�s\���B_eDj�J!�	���%|}�����3��}g��{����D�[���2"Z+��p�쐺���@�;�#?kD.��~��7���«:��O�S��'��2�N�{��G��+��A�K�kȦo����V���˛�y댴�3��E���MfL�)���T�&�����6EZ��]E��y�r�BNo|�_�6ZÂ!f�k��6��O�UQԀ!$pqCj���l���yɾ�Q���5(������I��E��3{���p��z�f9��%�7�u_����-vG�S&���dL��$9�����cu,L&~��4-F�*#n���e�;T%���C+�3$�g#�l�ps���Q�G9
+>5�:~EXQhJ��{|��B��T��Z���BI�WZhf�I�*�0?RҬR�y�1ڭL�$h.y�H"���}��L}�*�(T�`�8���Gk�+"`û��ﭥ5�����.-U֫C�1�vY\{��m��/9?v��$�[+�S� QS�����Uk�@#R�)�[qaa���'��CP���Y�mci�zse��#�^O�zݎ����8j�tLi�̗U�+'����a�����b.Ƥ�.k�
��J��,_���9�~�5I7����1�*oq`>7i�}/+u̞��{�'�u��`�?�7.(C��e�ӣ{���;"/��"ѸŖ�TQ�?��zmj�c�o�2����a�A��$	���M.�5�Ĥz@��
?	b���GH�Xvn�<���E����f~л�8�˷�g3gئD�˫O�+p�*���Y������׃߶,����:��?��'��>
�N���c��'��G���6c�P�-Wp���Tl�&}�ҧ���M[#S����>vIOqau��//���zd�v������m�^mد�*�_���d%�c��<x&��9��Eg�#7э�Ģj�,��/��I��y2TRO�O	��ϻe,E٤�j���
*��L�0ل��{�ڻl���]���|��^�6�H�<kVs�ǅ#.�(�T�c�o<`سAJ���Ũ���Ƙ!_{�4G�Z�d�u!\�Z}Ur��ۋ�����M"�,����}��ل�{�#�U�s�P����I�t�)�T�f����^k�Z��PM����b���R�UB�ؒ�Ok_����+M���o\x�Z����E�͌�I�g'��[[�h�e�R�>K��鵺���{��]W�����}N �Y��b��� �jT?n�ς����M�(�{���ʫ�?�XTe�����f�8�Ins�=m��>�?~A���)�i{ ����_d��m�O.��M�l��ɒ�)D