��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�&J�F�FOΙ{`�����Z�$R:)T�uE�3ahߵ��H����)!��������s���0l���N���G�F���:{1L���^�*����l�3�
�Zۭ���
q"�lν����sc��qI7w[wb��&�T&�`9q���.5!�:n��^F����k�\��쉿j���y4���,Qٓ��'eF����ը�D�ˤ�v�C����,j�I��8�V�\���5�^{�����?l,��>��M�-��3�,�L�h�}��l�����x�!)[~:����6����K�Y*٦� ���"�l²yh��&D+�ҟ�mc�M8�U3��`��J<��ԬFuM�j��&��	�n���vpX��(�Tܽ��AZ�9j�kg�1&[\l�$R~�a����1(�y��nA5eZ�ѧ�!� �;��"�t��.e#;��0�WSW��ڬuX��`	|�ye5�Y,4����H��F���f�w���ؑf)s�R�7��)���d8���I-蠍`y���\Ӯӱ���?н��� �X��c�=��2�q�8��:=��X�J�%�ͬq�DKg�qmL�	^���_�z���+i��>�M9)�
S߄���;Z�;�œBÐJ$eQ�)����h|1��jZ���D����y��E�I��W�w���:�Д/�zg�tĭ	Em烖 P/`n+p�_a���x��i�nm8���a3<
�F���J����1��K�_i�_��o���n9���.���k���9yQ����Z�ى�T�,�+�=��a��b�b������ `xN~�4�cbS;�� Q��[K#_52y�R��2�K^�P0�Yj�Y~��=����(����g[���3�h�IΤ[��bb]�jV��_�'�N�,���ϫ�{a�K��`��0a%��Yi2��/lX`A���c�O�'�^�'� 4O3)N3����0TH>pј��'Q�Tg"^op����ql�Pg�����hƯ��^ �E����}}��ݸ7�bL�R��\Lŋ%��_V�6 �B\�:qd:��8���y�P�,�a��K�A���}(p]h�3��k1�*�e��SuZ��sH, �n��3�0^��!�l�2c�g�_��ӎ��1���g�cF;U�?���pbWl@W���LO���d�n}sV����E��Gß\��i
v���«zqt�O榱`�[s�\7^����iG@�j�W\��F�MZ�hW�zDH��V�ޮJ/��2�u��5^'w�\=�	�;���!�u_;�f��IC6�!ݙ��(�(	z� �[# mAA;�5�j��?8)K[�[����%{��t*�XY2�-��ČU��%#b�w0$Qm�5����&����x�F�rEM���W%V�� ���:>=�i�b��f�B~��ADO'�Z�b��Vv��~l/#G�E�����"�6&'�n�j_>�K��<��߭�i��uB-	Ked�D^���l��l>�63;�����x1�ld�y
���U����$���CE�:��[[�Jt(��c@����vJH#��׈��&o��t�]����C�)�Z 3��#�&Jk�J�`M�U�)<�8���a;k�z��� �F�����G�o�-axL(��T�A�O6����-xj)8_��N�Cz&��Bv��o�R�낑c�����_΀���F$�nj,��蜶b
�������7
n�(hBQ���K����	'R�j�\Ӝ�ҫ%��WJB��<dPo�}fl�="���3��g�ځ:�"8�0�|h���Wh9@��!��a�ۦ��������J��U� E��2#�Z9ܙ���.��l��S�� ����e��5�^;N���y����C���R�U�n�d�m�u�
�i�,�y��!�[������4)�L�JK���h��F�+����;&
|-�O&��FQ{�w���x���b;Q���g�o��C|3v�z/��OD���[î%2�Q��q���o����T�62�ɚ|�o����c�k]኎�e�h��&�G��a�=�5������"T��U���}"�O�a������:�\��K�`�UBǸ��-�¡]�i|Äݶs�]�
6�{�۫�;��t���t��y��-��;q0>ɜb���<:R#������j��V�)%�pa�yN)Ť�<�Kzd�[��Lד��x�p� ��=b���Ԫ&١M�qc5GĞشZ�i���[b���2pJ.vy��}��<K�.L�Nd�+#6@�bg����R�:��!W}���{RtK��"]�F�75�7�����Pė��/Nz��ܱ�QkCTr�k[=O�d����QԈ�y���W5=��D�.��̗'W�rƵ�e����'iN���Z�"�iN��%|�奺��D�h�I��A��q�#��s�n����`�)���*����'T���p��q�fm�e\��k�Y�dʔ�P�~�
�@�g��v}�~�`R9���C0���-��ՠ>��˒�Dp��4�I���{�N6ы��܂͝�E��w�)��M���nj�Ko�Ea��z����sY�x�H2m�8� ���(� �r�CQf��A���6��P��O/q���m�7�7�ܠI�5z3q*8j�1X����*�j�`�:ְۏ������l�E�Tb刿�l��)�uML�;�*.��+�T���ү3��\���7kv���S+���Qx�Lb��9�f�&�$O�P��6���P��Qy��w�c��TYs�9f��yT���P�BFȟK�N(Bi�җ�gYy<�%����PT��@0}1��Ѐm0�� ��VM���Ή��o��j�+�n��эm��p�=N[hF9�¤^=���T�}$ �6z�M�i㼧�N��Hؚ���}>��".qF�3��zH`�x饠�����n%v[M�t1���ف,~R�7&.�U�t1����ׂn� �m��k5Z+�Ա}k̬!e4�F�).�����L86��g)���*\���8�Yn�s˲ťJ�9�+M�9�_1�V��gV��=굤�