��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ���v�$;��a�k"b���"����Ģtg})#P������Ӷ}azd	2vmư�s��MUm���B��]����0��3����Ng�s�_9Dm�$Y�҆s(�
@�C�1H�H�f%��ǂ�9�"��V�ϋ���Vpa��72�4�`4Ut���$ݭh�<s�ie#P0�
A �.���s��� ϶A?����Wޛ���M��#��hb�X^V���k��fG�m��4���Z���s�b�*`�|#Ҫ�;����(*h?��vo��*�+�'a2Nm�1?fRc��D��V�4�d�z��oҐ�Y��{�N��BǛѡ��6�$���2~#;��\TX���#�͊2����"�����|�p�uG6�;�&��|2W!։s�Ѻ)bRy��$�̛acv§�b��w@�)��͓�}6���* ��Ț�$��Ί�Tܥ��l�T2��kS�ƣ�
|Xg�w�jW�+yZ����V���D��<�<,��eBO�����\�v�<���ȴǈԔ�^Z�g�/��
�b��B��R��-'xFYڶt�*��A�k���,iU�_�b%���^QG<ߐ-\�yxa_g����U 辤ԡp�*��|e� &㥵��iΒW%BkA(G���z8:gߺO�!��<�F�������"�#�+�P�a�Q�h��r^���-��m����bɵ�"3��P�W'�0>P
�	q%�w�˿�:�n�&�&o��V\������Byu�L|u��CG}a�l<�	\7qr��N���w"a�Z.օjWo�&L:k0U[��%}�DvX��r8��7�a^��:�hK�:��SAAK�L22����f��
u����c+�ŰO���d�g֩GT��m�l�Oh�4Q4�v���i�~�rx@��_�黤J���U-�fӚI�K�40�G@�2����/ܹX!6ޓ��ɞ�0�����$N�o�Q�@��G���)s��}!�	b�2ѵ�C��pMXZ��+��&��R����q]b�?���M�/�x���Xj��>%D�~�Z�C��T#k�1#�����;b��Tee�1\
� (e'�=��͒j!K�/؟�����J����l.���,ﵵ��f�"�>]���n�N0+���5<����i}��f<��h��LYsFS��+3�'��6���i����H�]��%��W��ǩ�ѭY���5�rT�L�Y �z��pyV�nO����%7^uV��2�pJAx��\��6Iy���x����2w���m�5���#[��K�R+����1�5����{�A�Lz< g+&��I�G��h��H�����s�jn�d;;�*�ݜ�E��,�dU?e�%�:a�{���a�?�ޱI���H��ӗ>�	��������0q,"u%;3( ����QTx�zKm}�Wx�꓆89��Ae�MФU4��v�"��W�`�l<�/���5��(� z�埱�k7�!�~uM���� %q�=�dQ���e������q?���6��y��8��G�<Z��j8�gi�/�����O1�ώ@[.~��D�Tn�#�6�<�/�Tv�gѢ,k�X�؏ߙ^�`܍�)I�1/l�0�\�D�k���^o����w�����P��J�RYJ�3u"�9;�?�ѫ����q������s��_���c���O'�Rb � ݋�x�O/��g���j����"���� ��!���m�*�:���5�����e������0FX�C�R��D�Nm_��ta�k"��(�G3�r0�
)�Z�vF��9�y�d��~�Z�֖F��Ҩ�E�,C��gԺ~'UĂ�(�����Dm�f�R�k��ć�l�]va�tT�#\m�������L��W�!ui"�8�����aD�J��1ߕ`����n嵗��oO�z���Uo
�l����&�RQK��!���p�H���WN�� F����ǹ��4ta�is�w��;o^�@�wjzd9x(s���Q����I �.SJ!�?�W�X�[v'���&;LH���u�}>A7&)K`J�oIFS� ��)��L,�g��RN4�o��׳�;!n�d�`�>�t��c������&X8$��iu��U.����a<�	�\ 8Wc���g���r�__e/*���?{Q�V��>��y\>bB�?�oö<[���F���W��ֶ�E�Ԟ�z�'=p8N���Fʈ������C��R߱:*�֥dԨK��x��.���"I�S�zS]�S��9�9u�˘�/k-�qÅO?��]�j����MK��9A�Y�hx��p1��������Z3D�r�FG���)�?�5�e��vǟ��8�A��)|Ֆ�X@�a�G��2C�t5��3�_+���bT�2�z� <��,;�����l�jP�D���53!��D:��y�����.D7Ed�zX��G/D���C'C�J�i��}d�&�(�D�*����>N_U%��#�v�������'oX/�mT΃3�����(��O6D��0��ΊHz��[�'M�/�h��3!�m[��2v��6��<�L�pdڼ,0�3��j��e�
��{cq��0���
�nd
�6�1ޏ����_�����]��ԣ5�H�����8��| 1?#��[��/�R\&V�[�,J�y���T7Q��%��'b��T,�׋܊�P@�!Pz�WR�*mH+XA��D�D�Ѳa5���r�?{V���#c}��y�����^���:��B����3��/�gyt�؇��	�?���@�_���
0M�"�8;�3���߄��^�j�_Z����Ȩ��#N��q�����z�O�lПi8��Ȣ�B�r3�XT�3���.�8�I�̂%L#�q����th'�hٸ�\��@�Tێ�z�SH��Kj��7ʰ3�ySS)%�ySӓ�@h�A��z~u�܉�u�Ngk�t�	������7�حpo�TLV�Q���N���ܰ>Vߗ�K��4q/cɽk�Ђ�Ô|�����f�LT&��@���0Ӟh�(a09�5)����%�3�-H���r��Ӳ��>1M�<	��wpU'��%��G���ؼ-5Xb���6�lI�?�o�K9! ?�<1ו`!F�UBh�p����q�ւ�z$	o_�4�OPM.�v��*����Exd5#s\T�n�X�Dd_?,���+;�F�B�;���I���!^(�Dץ˧��Q]b�پ�E;����8���Y9���*��|:A"�jiE:m�`��m�*�����}h����p�3��.���ʢ{�b��l��q弝s��˄ ��v	SF��������|�u��FB�㗺��L�g�r�:���\V�iUV�}y+�0f�E����b'p���U���6wL�G{&�U?`�h�cvF]�@�3�J'����t�m^º"�}"B!:48�
�6"�oM,��|"*r0�R��xe@�1��j,ٰ�7�ǻ���Y�pu�s�z������]���z�>�3�N�S�@s|70;cQ[]��ch���7����m��Z�h��k��'�c�<bg*cN{��ᓝ1:���a� |q\_0 SZ� Y'p4��o=��1B8H�c~�zM� 7A�y	,K������ꁺѰ����6�v@��GT
9�U�o�R5��2)[�K+)�^��,�<'\U�:���:Ǝޫ�Xi�	%�nvѼ��g}�I��p`�w����kì{��j���
���M�ܬ�����}��U�Qc��]�ѻ�b��9ʧ~�5hK���I��Ѥ���Av����2w.��ĩe������ǬGׁS$�}}�+��uA����"#,̴;���ܜȿ��8-oS�T�IoV�BsH،w�ϭl#�� /�������wJ��ѫ�xD��7{Ik��������HOMB��=�NF@U���2��v� FB�'�,9D�5�b���ؖ�T�31�l]NDN��F��k`�m� ����y�w܂�=ed����7͐��5�h,�V'V�K
����B�@�6UO���mr}F�bn]��5%pjPT�~|h�^4_D�?��Ș��)�!��ϽMP}`Y��nP�{�r-�����������s�I��FIʢ�p� �x{q�.;~�n�'�z��������O>�4*����<����� =�n+z��[�fq(�1}��({I�	~>�� ����������v'��V���W��f�$+�K���6U_�l/�!���&�>n���H��I���o9;���xn���
r_��ܠk��U��ԈΞׄ��ҽ�9�!�B�8û��_1��o{�����-ϼ�z���4E�(��%+�}з��Y�?)��h���퇌څ�e��{��-?�������L����D���h�z��ν7��P���`C�c�+�'�t� �=N&�t�4��S���6�^��75r2���hu��wB�{~�&!8t��r���	��J�l/��K4�[Ӊ�J+C�[��1?]�*�,��|O~@?�H�ݥ�;� z��Ɂ�=l��a��,NS��U�c�T���CK�� ��ɺ�t�Ѣ���c��y���nM�JJ�md�녋z��[G�զ��%f	߭���F��n�����5�f �v�B;��ɵͥ1Wׯ�(���W������ Hy���	����V;3��W<O�9������q]��U"eևɑ���q*~�I��!�?,Ԧ�v�-;��
�b���Y���`�B�l 皞����@ �	�怚�3ZQ�0b
�^��.�"6��K/��0���B�a��� ��y,���їt�(�"}������Cޡ满8�!w�I��c�9�j(���-#�T�(�ɬ�6�Y����+
A�	���u��*��x�q9q��	CTպ��k̽!BF�tⵚ#V���qN]�$�dG8���8Q%
a�H�2wƗr�������vJ��*�#\�V���O����|o"x粠��/�./Τ헸�k�&���:�[S���6��N��V��%���k���	�0ݘ��U�23Fd86��0T&�ȷ����Yr��x��2�����sđ5�{6�p��C$�Z���Mx�9��62�o��Hʈ�������9�r(�x�5�=b��,�  o�9E�������e��$�{����r����Op���\ht"F�8"nF5�y����ҋ+�8����!)G)$����_D=�7k�����c�Y��Z����_q���ҵ��{r�Ѻbw\l͏ɒ��ZD	H�8]eIup8�2TL{_[g��.��MM�M+߹�f� d��Y�%�-�=U:Pp������W���k�Y�͎}Ћ��\o�g�DIET|
pNP���T�K86�^&��X�$�������;�O�i��񖳩"p���h_�
�H'��;>� ���v����qDPg����1�az ]a�S��I�7���z��P3�3��nݘ�K�8�Xe$(��#'o�*6(���cod
}����Q� �;�fn�w%��=�<��t�BY����0���Rv$s`�����N��z����5E��ݭ�LA���lY3��yE8^��e����w���$64u|�>�a�O �� w�+o�WdxYV�nb�N�T��r�z�g\[�p-�'�ߟ�6�֦�����~��e]�zflD��K��Y�ä�:҅EP0l�a�^R���b�&�j��1�*t��)�t�������C��#.�	���>8�W�[�)Y��}�-�vF���?����]�����<�J���D�}�s
*#�v�F���%��J�|ow�!�*��,+�X4J?3h�INs�Hn����f�w@��cV��$h@���+�(�>�k�����������
�TIɂةU@우��c����A4�@bS�7%lI��!���8��@������:&�xddd50��~���8���g4��1T3�~{&�8��H�Ęԃ�!0I��+�#���$�a]��e5u�^��$����~��'�P�W[���k��H��r�,����,��m��w� HSWU�#�U�B`��K��S�5S
�y5z�c�q�H��ƕI�z� �Ύ�! H�Bžh�Ŵ��:�9�֒��ǉk*���è��y��~t���V5Pw��f�����#	& X)
����u���������XX�菈o��F��=_����K�U2PQ��ǥ�)��'���Tg{�^��n���SEP��C�����M0�Ǒ��R��%����:��? ��P��7�b���U��ꕂoR��<m�$�X쪜���Uz����՛)�ۍ��4�\�Y��)��d���8�b��Ã��z֠:�Ys�p�������:'L�}$�D��.��M��o<���(��73�?q��>-�`e����aW!sˣ9o� f��^}�72�V$9]�񹛯�]�.92���z�ֹ/��jp���8���� ��i�ۦS��#P�hab���g�-���`�_{�'ab�.r�����H-��E�!~��b�4Y-��n�)�+�Oڿ��Q~[�W�Z6%W��ËY�0�5k�D�
�3z�x�W���J8�Ōw��# ����,��]���[�s �L�i�#P����v�(}w>�V8$�����I��_����<%n�
Q�Zҩ�;՟̴JȞ��L�\��9�{�2<FPo��;�Qg��l��+ׂ�UƟW���]��p�}������\�`?�Iǀ���gBdq���֝��ͷ�6?Ʈy�����6�	��I;���MHe%����<䤵�KD��326������ ���*���7ʹ�Tg�R�s��
ϫ�p�NzɈ���X��tӡ�[W�_�_<́�_�w��!�����$�6'��������l�%!��q��:m~�1��I�^z���^F*2��PG8V�yy%Ox���#��+����!�;�3����J��%��5�R�ٯ�7,�Kl;K�ܓ�����	Vb23���0j���!C�Uj�F�31~��ą�������Y�j����֓�A#V��U���<b ����^��{�b�{�fhX}mx�*x�xvD58��hQ�՘cZa��qϩ�IgH	I����E�-L!��S9�^��/e�O8\����_B�a��q]�����}pe�oe�����}��`��Ԏ�'�JS��R�hMm+[��������P�^52e˵�\r��wT��R�t�f+u';��#�j�m���)W�I࿁���x�7g��]�4�������-P�0��G�*�ߤ�����z[���W�M%����dӆG-��}�����-s��]��I�@�*p��}\ʢ"��U%Q�^.x˸ڵ��.]�*H�d�+��%��F��K
r����."�(r��1}����+�Qt@�c{�_��<6};ʤ���P�N�z*�����%V����6�����X��)1b܇c\��4~���6�	�Y�*�p?�����X�@� ������Z�s6X�" �����R��D��˧�@�7-�T�&��gQ���/Aة����#��Q�X����2��!�Iyw�˄����]&��\�>���Ո^���|�����u���u���4!��l>��h��A��k#з����xErh@��	r��R�����M������8\�	�E�T���}Θ�'���7%��j�>��Q݄3xq��/�F(K�ў��AUJ��ߟu�����ŀ� ���"����>i���Ul��x��k�N�=@t���z#��v3ɞ<��y�=X�)��$�wA��`/���*(�F�掁�6wz3��MK��r�lS�����^eK#��͠�ZQ]4ߧ����|�k+��憱����O�W�>�q��Z?��>vϠ?�K�?��vЕىo홰=��
"���s�0;��E>O>��8:%y}hG�{�Ft	�lʖ�� Jg�#�?� 8�`D��3Zu�0��WY5k	/�?�eA��a? !���@��[����Fv1 yu�F�=u���}QmU'�B ~>���Vp���v��waZ؁�B+�Eu(5�M(��b�7jse�av�򏅄��ݜ5eh�d|��'�0�
V<b{��	����/ׁ?�d���{���P~��%����<шM9}�B��*�� 'o6�N�[�uA��J6t�F��(�=�%���^z2��Eȧ0pv�̈#�v�"����V����S�I_�B�I+Z�͉㚥r.��bL�(�}����^��#�{��]�x�|��*@R��x����qۖ](�2�ӌ����L00��5���
+!�5��}����qY�C*�^��A�]��M_V�$wA�=�vĐ�܃�;��-�3y/P&ݱ��N��(5㐠hu�<����#�f�Ÿ��w]�������z����[�v�������o�~̐���S,;��+�|I����
غ�7��?v_��1��cF�G�+*2rW�v�M2�ώCL�`�|��[&ʝ}P�꽕):B�_��c�nϺ��V���N����I����{���i�a�����x})uL�/�F�词���:�?�h���ӿ �2�}�$���N�^������%�Y���P*��C���ߛ`d\��oyC-+�4�`<S?i��7��}߾��9���X�e����}�{O߆9$Nln�]=
C"�S��'�[�M���U�ʰĥh����Z/y�d�����n�ӂE:2	�Bn�,�����1;ˋ�y3I��N�J!L���uJiNR6E�[�7��p�kh��3��6�rZ&���Y��[9��g��@�P�^�8�"�.IpzG�c=�4E��¼X��!p���f��Əu��3�.�o�c
��&��b�XArp��?��}�к�x�;#
���n��1�Z�+}�k��[��T�S���L���锭XϠ����~=�h��;\�9R��o�<E��f�v��|�[����%���|
����T~N�gk�����NVYT9<�?�[8����7(k0��O��3����>J�r9�N��X�ؠ��=�+��W�k�����&��}1, Ŗa��t�� �B�J�h0��ǜ�݊	.J��2��K_�[�a./)�Umq�I��1�u!�Q91N��w�k!͛^%x�OV-x+xidim�E-��9#��yu�y�a3��]�o�zq�=B�D%&���.�<�}x���|Sа�&
-��߃�N���X)�gR,�g�3%�'���^GF��d�6��� �#�J�]��@p��>LZ�Q���_�2�%-ݸcSS�đ�����0�M���=��fyR��gy* �8!�Ě@��\�њ�����?�t���U[e2b�"�]��斫0Z��sn��K=�*��f���fxv|]�ӭ����=ۓ+�*�j˫�	�#\xףh�`Dm��U���l�P���MX{����9���*@�������-3H_43FCd���xõR�«R	^�`})�<�� 4�L�q��uPa�l��6��
��:]:c�	%��N��">��W\V���׼��n��O�T_ϡ���<2���5��=��-;�V�P�A�X�ѥ�45������jB�bę�i坯�t��U㈀��zA�-�����[:�5��m�p�(�n��>��:=�6��$�G�Y�D� N��e���}!�q,5�cL_��%�4^�Vč��Z}R��c�T6�P�48Z�7ˢl��X�!�s6�B�摫��t-~�P�������9�sT|�0B���10��e��=�#B����P�,�v� ��?�Zd;�	5��פC����ϱ��[������!��H�"{���z�i�0~�Q�ᖪʂ�$��>As*���Ӎ' �I4��L:z�g��]!+�-���K\tU>O��vQl�5�N�8�����,:��%��2�}�\��#5� *�c��e�+�nbD�O�R��$�RZ��R�E�U�R���(��r]����>j�M�L�+J��-��&{!�UOh���w�Pk�Ҏ5��ҦХZ�Ʉ�m���o%Z�4q��Z�B���j��%
Ėh*�7u�#�b�Z-G�2�Z��8V������L^�]'��o��od���O����K0#�ݻJ`���g�ua=��M�.���ʺ�s:�0��}eU�Rl�F*�m̰A�B1y��������c` �o��2O)c�@��֕�P�%@7<�8d8I��'�Ր��A��S�}��Y=V �ԃ{.��@r8b��"�WIkrϖX!����u�C��O<5Ii+X˰���ɭ���qnم'^���ȟ��c��c�IMmƗm��f��wQ���@�0I'����oF���u�Y�b�}�s��D���ё�u�4��V�m���Fl4ʄBT�D�E�mCQw�
�e��&�"�4��ǻ3��M�F�Y+�ܹ������Ukt�5�7�>y�8e����q�l����`V�N$�6e?w�� g؃6��duN����J#�$�� ��	�Mz���Oee��/b�U�H����=���R���<�T(r��V�p�i�~䢉�E{R��MҲ��t������P+`�ORr���!��v���Q�;�O-[�Z����ޓ���<�� �+5)���xlI����w�ym��j��xB �p�r]J?A��Wrˋ��}j�g҈�韘������<���R`n$�˻�JF=��S��1�g��1��/��X$`X�BDD[�a�ƭ����1�%!�c�9+����̪O��zs�7�M��'��ImY��l����m����ɚH�v�yL�4?'�Z��x������5Bm7�B����q_��;Œ�q�|6rJ��5r��m	�&�����}!�Rs�zh �Cp,Q��ߢp�����#增-�r�/|O����^�q�y����F�T5JGW@m�����L����P��U����%Q��~+���>��� ��{�|�X�×`�,�2C����	6��ǚw���$�1^_.� �샼��E�L��{g �gn���,�Q�%n=���Z]�+ܑ�l糦푟���x��X(���Ω��[ʍ�)�^����U�|�<Nn����,w�mx>sV�~�y�`Pǒ�5Z�,�D�_���pz
�F�<ؒ�{����#\�B�UO�=Φ��GT��8��I����͆�Z]B�f�E��1b@�������y֩���aX5�;���k�u��x��B����b�����AO���4>�TG�qaȻl$<(�u��@�E��+|6�R=��s�ʆ�
B��n-��Ǽ��y�J���GCF"���>?�(��,���~°Se�,�����c/kC�e�r;�=���
,�?,�C��0l4$?��-�N�C'2��7
��g���u��z�];����e�!TY���*v@ �E��P���'�?_$�����7i�j���T�7��G�T�� y�#�D��.uW��ȗ�U�t�ڕ/����XLSI��Z!B�,O�FQ#����dRw��e>P�8s�����O�Z�l������8��f��T�q���.���B���
r��A�����C?h�
�Oe�6A�h��V�{�i�"fi����qIs{�(��/�oʅ`xմ*y���շ��#d��sƐ���_�O9��Q[�X)����Q�Xf�o]2����40s
C���"�t�P�B0�vK���m��ۊ� ��A��"�W�~{�5ֵ��z�Ьz����eMy|7��N��N�u��?�׊��&(5�V����ʈ"�P�$�_�Ejdv��&�[��ہ��; ��9(�.��ݧ�m�R��8/V��ə��A������?&��;0"{n�e*Ya9��L~~�F/�V��V鷭!��nCo��]�e9Ў,��~�{���� ��o��@���SPlW8F>�ʻEY�87��^�:���UY"j{2�A�|:ҥM�C�&$j���+:�(�I��hHz���԰����F��� �ၮ����r��b�g�[�-sa�ö3��Q̻F���#@�J���A����k�wI���{v��F�8G|��C)�P쵀�M�t�+����n�Ʊ�Z�JA�o`Ȑ)�-r�f+M������?��q�vFм��b���c�#�pϋ�~��=�ZQ�H���l�Կ�6�s�/�u|P�)M_�ЏRf��m��!��e]�g7��'��"�/cAr���+.�8�`��v��M�2���[�����|��yV��݃g��':�g�ޫ�S�Bⴣw�g칻�"�=���F��f̑>�
�b�+�D���z4E�3��1�0s�	��-_��O��Sx���D���>8.f���~�ɓ�z�WZ@���u)"���]����?p4��t�y��c40�Z��,?J��=f==��@m�ȟ��j�ߦV����eK ޡT�ؾ�(HQ��2��"��Lฏ��0`64M�r}���
M3nA����sU�.1�z����O)p����-z�a<��y\���s+���=ʣ���;r�b��<����6,#~�'�,�0C𢶄�㛋q���IE�@x2R�Cǆ�n-g_�T.��+�*�Y�%�r������u�����C�'\�ґ�yP�goV�^	�N��*�&�8[mu@�`��)v���e��!�#�*˓C�6n�\}�'2��:e��+�`+!g��#�Y>