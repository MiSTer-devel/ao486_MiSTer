��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չt�-���{�\q�e���	�jE���B��N߽d����y#Y� �*;=��4���k d%e�A����g���]�-��C'�I"vHjF�ʍ�9B���n�Nƹ�5z�0<gj��M 0�9��"��ʳ�\��U���W����a���c�I���Q`
��(���[�ܰ�<t80D�������ܟh
8��4%ZE4�)�x��T�\���ٔ��/(�ewP@I��ߏi{��(�b��e(7�	6�1�kRl?>L�s�.}䚲���O����;��P�@���
A ġ�7��g� ���� ��8�h�|���+��JJ7����=�
KQ`u_��[�Ԍ�ԗ`�;�1e�=��C_>c^g�{�F2�]��x���\!/��f��N���uۄ9%*���_��.��Q��*A��0Y�m���Y
�D�v5�a:
 p��1�z�U�1��V���,��,� :�>W��ȿ���u%wx�9��ɄR�0�lﰠ'�Q�ȑ_�(U�Q��&z�	��߻n�yc�&Ԉ)�T�_̸�Z_�()YO�ή�:�� PC�JXe�҆�P�=u��Z��Q���t�
��n�~0���4*M)���
��>}��S+�D��@G��:���W�a*��`�^%�(�\�l��!&$��G�mړ�׳y�7���ā��R�a[Tl�OUS�OB�؍u=� Y��b���+P"�U���;G�^�'�ܷ�Ix�T+�q��2oG���]mH?�*mƔ�J�BgR!�-�+%��lQ^�|`�9S�
�U����Ч�6��&sd��5�X}����:�$�@+C���g#�dZr��m��|L{'����?�8C�v0]��༞��?'��/�!j"�U�����
�5�J��6R:e���$�&~�"|MN-��SV�`U���ט�t���R�e��d�ଭŠGn 
_,���SM`��!; �AZ�صUo5@a�Kej��Tа1)���X�X8���$�/z#�������"��X�b+SF�yTz{&ͽ��w=N�Pyo{�*�la"�s�m�8O�T
eؘ�ea߄�岛Cg�T�����B|0/�Z�flܜ��y�O�8h�P	ҏ13�+򏨌�N��m}��4C� ��t8��$;w�Ѻ�U�f2)��2�R��:9��yJ{�	"��7��q�h\HĶu����QzFUXR<O���d�	�M�BR)�w'r����Mu�DC�s��x~Sޝ�K=�=�ξ�ȯZf-�s��律P͡�2�����9�����ȗ'�B�*�FQ!d(�K� �D��e܍�uf+�q�f6R�:�w���������P�#��I����_�lԁ��E��X�Xv3��{%�;����t�}zP�n��'�"�5���gs��[�mD����ᅤ��/L6Yy���* �m�I�|�������Y%;�)���w�e�x^�9Oԟ9�<xa.��A-]�|%�=b&� �X�{��5�dpV.D�������:\���ZQ��/ö��y�g(��Zq"�b ��r�ܒA��6����d1M�p&^�D��q^h˵׼$9r^�������