��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�]��G���fy�����EEP9v�.����(��kL�|�uz��M�D�=H���4�tl|��M�����?�������p�&�dY��
Z{W�,zN������%��vvI��dB(#�6�)�Y�����eY�`���pE��O�cX?� ���rZET
:�s���L$��/�W���+��FB��M�nbB�v�,�y��U�{�OB�� e�8���Z�]�q�o�Ո,����<�a����ov��B�ɛ��BMK��1sL��^�`u�	�A���-�k>�nO �ۇ"x3�{��Ҡ��zp�U�F�t�.+�ɀSǙ��D�����u%Q�[�fi]���n|(�gE$�Ę�A%$�3�!�:/���Tm�>�B��F������#/�+䐱�wA�q�a#KW9�>��-��n�i�3��0��`��|��1L�����L�����<�qpp~����J�r����LA�:�f�mB@��Ihا2�U�7��#���$��Ƚϸ�~[�J�ؠ�_�SD��jEKR��u;Z��1?�c(���]�����]�`D��P���u��D�M��&7F�zD�F=�Ʒ(���M�S����ޒ;N+ �<iȥ�j~M��$��,�}���e�����-�;`��K*��E��d��_4,u$َa����<�-��ޘ��0&)��GbR��+E�Co/���cf�&33+��V>#�7Q_�:�O��}p˥��`9��*o[,9��%Y$��?�D��1C�j�ׅ��d�����ۉ�����RW$��MZp�^g��E�tT���q��>�-V�VW$M���7�[Xs9Orj�@%�|vn%"�`.s�<]*������C9)q�Lͷ�C��Y�ީg'�p'�#��O#!#=AİU~(�Ā�3�sP`/v�]�昻��'�ѳ����<0��Y|K��B1�ɧ>��KI�$�9ɳ��򛯥$2I�/{�l��w��RY�	f/���Aj�#�C��r�8�_lL�R�W˨�5��l���p3���t.Cz��X� 3Ҿx�4���Y� LM��O�~FzF?�Q�<�3�zo�I<��mZ*��/g��!c ��M��FK(��Nq4u� e(z��1q�S��G]�%IX$�D���v�no�J�-�1goC������n�/�$ﲎr��WK=,��PX4ϴ-2��4�H�]3��ڥ���3z��lɯH�(�5�M�����7�uķ�|K��u/:�iS7�Lo:��6V��J�T�vr3�"pB��BL�D�#�ㆄJ���~r}��Q0eN5�yQJ�UmH˥����4:&K,\�᫒rO�679��׋�?�3�(��~��5Rsem���z�'/�f��IH�0Zo,|�H�� �>��5�q�|�Qא$*2o��H=����<؋����?�۹ ZR�.�E�*�aȓ���_j�c�~�:比�< :���R&���i^��&
c�\����_��A\fJ�j)��ѳ��l2����(�[7a�>*y��j���u/R27Y�Z�xݔ�m\�p����(&̡*�h�����R��H!D�s���f��ˇ������`�f�?/��\�)��i��r*`�TF:R�aúˌ@e\�u�ŏ��}���Ƴ�c���4�k���GV*�/%�M3�_���W���S�\l�ȩ�"}#�'�k�`�>���;v�����1�TO�~����H�F��0�X�-l{#�-���E���l���L��Z�_m���.S��hȌ�OAI�u�&S0A��k?r��So}Y|m>�*��&�6rD�5y2�iƣ&�	liͥ�tŔEB	-q����$�mh8^�ݯѾ�}'�m�Ut(adbQ��44m������"��5�A�b��03�7Z�u�u"�����g'�S���vyG�<�Ђ�GJ� 6w�KOӈ����i��h����<Xu��M�0������焢?�
�y8�7���A����g·q)���8����s��g�Q&����k���p�%_$��J��OI���
��*ypI���M�����!�OF���{X�q?��e�JO�T% ����í�����@{�մa,go7m^��c����΢���շw��|����'�.��F3���u.�>c��r���-���~3���[t>�Ll��=r�l�� `,��X?�^z�Ϫ�N�^�E�I, �X��q���df��hH������lR�7t��*�w����;^{|��	G�ԧ�t�5X �]ؓ��~�E��Y�S�|�u����4����L�Y��r�?!2���v�G�n��ֹWբ��Q����	R�",X�عɣ8`׻���j%j&�ө��a��F+bTe5�T���jP���BM�v���"-lN�헫�N�$�p���,�a��Ά�,S�ͫ22�C��#"�l�z���L��y�d#�	ƉbwZ��7��&#u�bS��x��$�H�xym�>����@rJ{k(A���$�|���.�]9�Fu;���2�5�q��e�U���9�N�kWa�� +�&��5}����6ru
6�Y�F��p�&����$.jh��W-�#�%b%����=/����y�ʊ/�sp��[i3���O���I�	�U@of&K��x���-'��l~ �(���ܧ��7Ư�'%I�����Af�'F��y7�T'#��'>o$���ǴG�+�93'�d5��ڪ� �B��gj�z��.s=M�c��4�a�/�G�8�I��٢lE��Q^=��rS��XCXT蠭���3�Um�_���@��k�x��/���`XM�aı$�2ۖ�u�S�%����>C�lU�ؤG�OHcAON]�-~ʸl�d�C�H���j5�3ߓ	����ԖaS7��E��:R\2x��ud��92�g�O���
C��`Z��ǥܮH�����``!���g���r����UۙmG�q�3[ћ�6&��U~�>�D� �Z�b�wD�W���D곽+n��|�f�[����4UM�ܦ��!��^(C�
������&+��;����W�7?���1��ǚ�m=|e���R�N�>x�"�A��M\ˌ:��G{ͼ�#�|�Vh�Ӿ��٨��lE��B��HU������~�&�N��/}�K;Mw�u���[�H�wff�
���2El/m��ԞP�W���fֈ%"|L��ѐ�',�Ik�����J��m,CG�������e��1����@x�?@R\v)�WË�x̓�әFC;%lcax��+�d���V� ^�ա_�>��K<h�fP��Cce�Zæ�"W&�RW�:��jlH�M�V�iNڳDưaPE�s� y|a��9XƋ�v��˫ݘ��.T��3J����xQ6����(�Nӓ �����H�3�yێ`͵��Q5�?J�H�����A>��,��[Hu,����V6A���*X��a5�	�m�X��M[Ǎ��xk}$��e���q�b�ݽg�i��y��j�B? G�`_F-G��oL3� <PuM�ܾ�Ȼ�}ݩ���Ϩ�୚S�q9>�l�`�ͷ��&~4��Q��LR��1�9�Y���޶��(Ax�f�ֵ4h�þ�b��*�!�֥ʠ�Y��j��8%?C� ��s�I���f�-猂u���U���/�U��d���;���C�J��p��o;� O1��:HF+�X�}OԎ??2vm�{L�j�dg�S�)���(W�*�U�b��?]kJ"�Zͨ ��5��\�"�zZ����b�5t���mN�y^
��"���8�����c/Kχ�y��M�U�)�X�p��W��N-5e�P�ؐ��k��9|�^�Zϓ��$ǀ��A�=D����Nxݩ�:w��y-�o���v�}�F��_��`\�b��W|�n��Z���jz����51���5�#V>Xz�l��n���C��?��^��s���^��2حOĮ��Np1{�!�6�اLq�@�H^1����D��X�������ޣ&b2wx�������I��rh��V+����QC�E�=ע���.��}X�!�w��I�3����ӱW��>S�w�28�M��H�b���*�P;���˫�嶓�s9`���������e��D_��g�ߜ��Ϧ���6 �S��ϓ�Ѽ߇q��m6��2@ÈI�`U��wx=��^����|`�}�e�Yv�8T�������