��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ���� ���^S]z֬gB���<�O5�Gn��R�s1������g;׷��|���z*l�P�L$ ���J�C2L?�����N������1��2�=���2�>����PM!�GJK"��%M�nx�@�g�����H����5�HiuMi
�j�L������+xZ�Gew��u�\��c�J.S���W�-�ٲ����gCm�.�44'<$3sg��t�������u��ZU(�ޛy�ӏ$��\7��K�8Rht�>�;�X�c %Z���a�q(�r��A�:����=� ��~)jDMZ�|�y���maZ���.5�'�!�ۺ��e)�
��ә'>ꨚЖ'e$�����:,Y��w��ϵ0\�H��ړ�C6�A4ub
����\�Bs Ӏ��Bn��Tkƣ��UQ7Pr��n�-lk�՘��Y�=Uګ�e�t�1d��+��T�m�4I�2��xkF4b��|�'�f��Il���N����o�,�pc�y~��r��x3�����'0���!�����Lg�}=�6	����~����_b.�b�ų$���#گ��YG�����]��=�.B��u2K�y�o����>���o�y��Q��M��UV�ѻ��z�-��C������|O�!.m���aU5!�c�$/QRʹ���_V���A@z�ʬ�].~��7��-@̽:f�r:������*�1%�h���|:ym�K9�]������t�