��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��ՉR��6�b'����0s����_9��F��h�'n�����H�:�f[�$NL�̴R���K����`��8���Ɗ!�b��qQ�5���J�+j><�>��yM�A��K�}L�^>>� ��Jb"XuA�r���㣭��"v���@�����X���^h�n�L�k:Z�{!���G�0D���l}�0����,�t.ߦv��i-��Z@����n)�j���������D��3����V(|�%��$�ck�WkF#���[/��_��
�A-��֔��f�\Z�Zr��}������Q=X嶨ȡ�t �Ya��h)b�,�>��o��� �N!B{�=��Ԧ��6cβZ{>6g���!��}��vlg�uS�o�Dч��8L�aW((������� ��%��7�+E]����A1�~���� �è��d���2�r=�4ܤ�P��o�<�歏��h���chn���L�D�ԃ�x,���~���s�@E`(;�!p��,L���TC;��b�n�2�#�rE$���!�{Ȗ�D�;{�H�F�|���IX�A4�v��׾." !y�N�*Xs�(���`�?��������j��!�!����x���F��W2F������b��A��zB�d%(l���d�,t��H�)������h���@gӎ� �!�*�cz"xL�#B3����ב�;��ʀ��bN�ce	�=ڹ9�xf�$s+�YK(�K��y\(A��Ǜ��G�' ��]xf�b�u��:F��z����i(���DX��'�Ҩba��Q�g@�#����ʆ&*̭�:sّ#S������&�¡K��{{`�0�B�*6�G�@mK������Qųk��qA���k�����9k���q�'��x�ڕ��Č�@o�4�?J�4�N��_�fjjv�̈́�^�ʀ46nuY%]ĥ���4r�"��6N��8�0���	��+|�5k��;돡y��:��C�C�h�����'���K�U��䒜�2@�;$~����sb͜��;�/:�k��URT�ˋ�)���gQk+��9d�=�O�Li�z��,���f������>�F��0��!C�p�x�������bna�1L8�ϖ����/��і��.ձ��Q�p��Fv���-AE⇾V|��1�.�'�Fc�r󐤫wƃOerP��Fsx{�-,?0��٤�	����^�_�,����v�){vݕ3�d�Ŕ��ohqY�s���>�:�
�����[���	���^�f�~�A� ���?e	P&�^(?C�.�	(~���R�ڭ���zs��켈�yφq�jOT8Fj���*,X/(�����!z�O�OT��x�SW�G�G������1��AX�`2VN&�ʴ|���2���Gq�:�
XՃ�U��]ǞNNFNi೻hb�X�5��	2G�y����S�e;���h�.�F�q�R(&���M�