��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��ՉN�*�s�/a�(,�ʫjV�i�g�R�Sm��M��R��sS$oǦp�&��oE�M���qSش�*�M8%�Bb0�aAA�!I4(�<3����$݆F�UK������Gs:�'�ȋ�:�hO:�.�V�v��%�P�;�� kd#,���K�I�*�2~����d���z�]@����}}ޤ~�|9�e|�x(،CC�q��8�9%A��FF������9��N�+?{o��Y�F�Ɂ�[ĭ��)؍���G�mZ���]����a��b�v�m~��
���غ�;��P��6�U����=9D�,��+b�sk���>o؉rλ�ta�l��.�. w�
c���/��?���;���QO�I	x���$�+Sx�K��-��-˄��dG��@��9��C	�jS�^��q��V�bk3a0��P�ә�a$ &�N���"M$p���=e�>4