��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ���v�#��#�K�td�~th^ f~�~f��<�*��O[=�^��E��"�n���m�
ص��~6*�����M+S�2��YGݞU���V&	Wk*P梙X��xÏ�8J��ka�	r����~�hM�o�� 5���.ӝ�w��/$�t�T_l���T�����C��Z�e���%�ɲ�k�^A`��קR��<��|���/ ���Ҏ�(�.d9i.9�:P�m&�7N�����
)��ǝF0V�^��_�k�����y��$�jW� ����/u����,�t+��bma,幆�*J	����0�.��G^Kw�R��|hvx;3��:�����J���%��(y3bt�/A�|p�p\x*8��}F��]�Ns*X�o�-�����]�P����[�	&�诋xQ� y�����h6hېcM���bs�p:|{����ɔ.<O��EZ9��1��I��X{�F-��~�~Lu�4������_�Z�,�Ԣ�q�n�H|�T�I�'$�,�� �o�/U�V�������~A$zlq�U�}�@6g�]��s�%3��#k�O�~��$��s~�[����5U���>�=(�D2��~+��%�2s	��.+����Qm�v	�A;�'贱��Ouȅ�w1���,3�J��i+��=�f��0���:��^�w��u���xP9(�e�@� �H�%�ȝ�N�M�*�.�q������}T𷬒�C�!�q��YMڮVB���n>֥�RqN�<������F^و��9y'��ސ�";�n���e��k8��"�ؘ�%�鹿$���>���=�Lȉt����Ѿ%�?%� �Hҭ���2��
��1����E }��ݤ��G�$lN��'�W�!`o��_�(_y�'���d��)I�8���۹P1@�-��� '+qJK�{��%�<��؃
p�|ODfkG[�?zD��t���V�����E����G�e����x�d���0l�#R=�B��\e�T�0eO,<���&mV��"�{���,���8fӏE��j���xN&3��\�V�Ϸ�	���h��Drҙ�S=x:���U[];�R�4y��R��쉼v�J���Ád���$���{r�|�ǩ�y����KW����g�6�{�A�PS=b	@�$}�C��ZEJ3>n)��]����~2���Y9�4|�Ix������=��{y�Ǥ�g�v�ƚ��P	�S��*}���� ��Y;��0�+��s=F`P+�T*�Nq���wdWhD2��g�nƕ�;߰`� �NF�s�:��W�C|��j�E�A�ۿ�R������Ñ���	�p��c�`�Q|�-hꩭ�a���o�2�