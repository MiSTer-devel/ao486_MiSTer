��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ����Kq���V�C,����x�,�EZ�0�@���9�3�Ż2Nl��<��<�*�Y�s8+ t�q��M�a-�!Osv�y����HwztU���s%����P��r�L 񆸨Lk�쑞B���٬��͌���U�5 RA�u���#b8)C͠V��?|�3v�X"�R��V�������rݢ�#�gs�
`S���XTf�^fi�[��L�����x]���)@Y����cL,|l�e���?��i@�����"�*�Eg�dA��8UX�:)z��
D�pF�m��0��u���:M�C�/1���(x�3�I6W[jB�H_�������) ���c������x5����g�7CgND����d��!��7H�U9�	�rٵK(�<B�xd9�W�~����*�ݏv�2���O����W�L���Xg�v}/uU� ��Z��pz�l��
����ph����!*%}�
�X�R5`��Y�U�cOw����/*��� a�́"4����z:�ݨ����a��>����*�Qd�t��S�X0�o�̟pWh	Z�S����-�X�b�UVV�1�r�<�}���5!i�@�ny��c8�\,E�A5~q��mq��n)hy�]�'�fص]�T�D�������i���dw0(�A�a�cz}��[W��������2��Ԑ�】�J�"*��Y���t���q�>�P��z�4�ﶬ�sԘ��!�/޽��RD�	e�1��a��Nae�W~�����`|�4(w��fN�Yd�^��������,�n�8@9��A��l���&U���44��I8���'Q|yC���*>H������?@e���W�`��T�ͯt8`^�����R�b%��ƍ<�OO!�b~�ҙ�`��-��q�O?�ϪdL.��J|��\�w�gusqJ�H�vJ�Q��A�-(`�UfB=�*3�I�H���1�_ǫ���s�!����������˾�X:��/o��<�7ڞBa��\�Dbo
SHN�5�d�A|Ph�'��i���1�I�9�F��N��0�T�z���&�W�h����P�S8��x��fi�XZm-Jg�ɥ,���9�yN\4���k�
ë�2��z�E3֑�#&��z�Ws�Tl0�CƯlF���ε�k�/�0IЃCZ��%k�@����s�5���r�r��0m2�'��|H��^^6���h[��y�76���	�*�Z+@��ʘTARN��u����d�V����IZ�T��u5�X������v�)Pu�\���b�)�?�y�=3\{ZSԖyͲM���l8�3�t����0��.w�<�t��Ӫ�h0/���Ñ��� w�h1��n�=��?ő�+J��b�0f�m?��"�-��m0����Mt�r��ʦFp����F����pUt����Yi4j�(�N>Q��y�?$R0fN���?���%��f���[�X�x�9I�ĳ���7�4c���O���~���0rsl���(�u��n���U��BEz��9((!yޚe>C�PVZ~2� 	Mat�Lu��$������P�yt�=�XQ��
�v��bb�Y��Rn������~ >�V���ͭ]�g�V]��+|=�C�z�O"�)�!J?]�K�,�F��T�0,��ړν#����S�:���T�}i5�ity��'��b�N5������B��IR�F����X�Br����7��o��dv�K�X�j�<�_���
1B����4�n��8����ɛ�t��<����nh�?r�~�����%�;?G��ݒ=M7�8R} il��(m�]�:1|��y�z���W ��,gF�@ƨ����y�(��Q�����2��{}dT��]O���<��u��$�m��)�%�Nk��YܪZ��p~ �����X��s1넅.)1+Fm�1��r�k<�K�l����T �V��E��\����LT� ����H3>��n�>ګ�S3�A�&�H�w��o=4*���O[��OgV%����C푤��WHe^{Ti!�O�.fG�?�������Z��/g�I^M N�%˄C9�[6J��+�w$@��[7Z�Pi�<cx�\£f[4Y�ޱ�*
��V��N(͠�Πkr)���u?-��{zX^��`�I�*1k���?���B�G�a�=v��5������\����VH�:%�q�k��/l�6�[8� ����P	Є�&j�����'�KU�ih�t�,�v�jS�n`	�)Ѭ��<K��[�4�S%��˕$oL���A�*CZ�Q�����S�����Z��� H�G8'9�Tby�`rٹa�
�6�%ns��K9�3���~5�XV�6�)H}�ʴ��딌��a����4�R���g�X��:���ז,:*�x%�/uW�4N�p�=�*ܬ�F��f$CV��ʤ~���a����Ƣ��{��c��K �/RK�v�<n��Mc��5 ������}J� ݡ(N"������
����k\#΁/�[�1�4�W�.��J�A%��*w�_q�)�L�c�/U��W��1�ˠ����Qp��o6W��ɶNU����]���,�L�E<
k�LW�P�%�1U���E�d��p>/�����$5^ i\��A�����-��cSy��.(q�<��<�HOZ�'iYX��!QĘ�;�׳�0\'�ɔ`�U�FC�_1iAh����Jů전��F��57�b�J'L�[��[�e�Ϯ`s7�e��~�	.�M�����"Xq�z��TX�a��JX�4o�<�9�� �1V��L��C�X��a����o�D����B��P�3XC���R4e_;D��Cc,�j���P�&��F1�3��?H^�8�� ��`B�@�y*����!|+���Г�#��
L���:�׮P0��eqk�O)) YN�������|�.�_����z=�*H��H�!��  �p\��O�>5S��mW�0P����Է��L��\����S<F�t(��u�-I�]F"��i"(����b�Z��V�����{J��������|!;y�ɸ����1eOp'����$!�r�:�<evK���՚N��,�3؛�3�m�ez6D��3�r@����B%���rՉ�Y�xǩ0�N��e���p�������⃈�<�9{�w�>Is6�f|d�S>�[��AߌY����&��C��x�l�.x�`��	�R��Y�R?y�+]B Q�IvP���T'���\�P�5�i7�%���*�o�MA����:���U��C�A�������m'�v�[�XcOrM��k�w��i�QyU�����H�X{�z|K#ՠ��*e�+�ޗ[:g�^2�8�¤���	��j��rt���RD1�P��$�?�J~�H33(&��x5�����!b@V�e"��f��,Q@f��jRP�vz�*�2��,�7���3���=��l�1�$�8��*�7{p�)S��C�:gZ���Sp�p^S��Ov��%��E��l�.���Jz���p#�4V�ayz��*i6��F�?i���A
d�ɿ���"Ta�O~�@���Kg"O�'����1 Nˇ�H�DH��\3�V��wf�JƭQ)�s/2�{1ty����%W�����}�-�X'�z��&L�����+s5���(Y���o:͒�b���US!��G+�!_o��Ϛ�
����jM)t9Kt�ޛuE���R�� G!�����|e���X꨽���l}�oF웃�ݘ)-{j/�(�����%0�O���I���O��bb?��ܓc[t����B��A�)���Pf�%�l;.��Ǻ4y��Aɝ�� �� ����]�E�������Xz��MdP��A��.��$�ؕ{G�e	ڣѺ�k�e�mݢ���թ���".P�Tل�\���#c�nH��J-(�SkRs_P��pEvHV�H.��ڻ�mٲ���V#��R�;Sgj��c�
�5A	L��
��w��XQ�e���p�w��ҙ�PB��]�Lj�$�([R|V���