��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ���v��|���#��Ŧ������Nr�H�qf��"���d�8��ִl��� Lyǳ�U�Ԑ����?(��	����`�?}���4H**Y�U���Y���u��s���,7������g�LS?�+��0ZB�Ks=��'<�B��+c�Ϳ<��5}�� Qn�Iy�@oL�J�?�8M��w�A��l_��-h�еb�+�Q�y�Fl���Ѹ��j'�\����pbO��� ��ksQǚ�&~���jt ��SR��0_l�h;�S�I����NK�+Y�o��;�2,;~/*�V?eڒ`�ZA5�8{B�>9}��&�x�I�\~3�ky]�{��{����Eؤo|=,�m��Mn��Y�4W�]x`�$/�a]:Ͱ��z-�?9>בK��n�Ƕf�/�m�mp���+,�f���p%E(���Ql8���g����F���l�G�o-]��q��u"<��}Q�Q~]���ǅ�e�wF��V�'Q��1zHO�omś�%u�~��nTة%@SKiX�^킗�6����A��S#��A����
UB�tw�#Z��-K���S\P��՚_�Eo�=a��a�U��]N~ާ�@����k�<g���&S�W��F`�hW���T>����7�/U�� ��P�d�h��r��C�鲲l�j&�,�`�0:>���g-Bt%@�b��0����m��H���3m��s�����;����❢����t�4�8�z�ް�XFh�����'^0�jw&�^r40�ģ����i�@y�ѽ�vU�%�6>0c,�U�}�!��{�1�4P~�A�2]�ƶ���\�'�YyRw����>P)Ӝu��3ށ����vM��5$�g�UT7o�Q��h�ez�K$�|����F+00Qf�B�>Fӓ�=�2y��w`��n�q��
����Bq%t�^z�Ğ�ɜ��B�y�۱�oS<4�?|� ���Y�_��+1��-���\gG��.:�&����K���R�4�8X�w~.S�����r�񄣊_�Jщ�ɂ"���C+�e��urRV:�~x,��ɑJDw�2U�+7��N�v	�\���%
�h����cs�R(q	����-w�Rg���TL5a�t��$֪pXTI�Zɹ��_�p)���f�����jv5��&�V����8�a;!��Db�Sx������.�m~#W����K�&Ny��>�ܜ�H9����%������M9�����&��j��66���m2f��΂���pm񅂹E$�w��T7R�ŝ�;-TN\�	}Z���D�ޖV�KmJ���V�y�˾��	�ݖa*`��j;���9�vSRl��tV�)"��yD����K�����@�ⅆwRD�a4x��ĩ��y3f�z�������=;дt ���ᐨw�ʙ���>�a� ̿�kw5q�Q�N+6�g4�H�&�����ƒv��J2 %����8�x��6�:'�꼠w0�lM�_�9�
��{��c�Q�m�D�Dbr33������e�N��U�Y|�.`^��{
��"���n��梅�0�����P麿[����0jQ3��3t0�"M:e�m�`$���Y���R��Y��YB�m{�M5J�����$25'a*����� ��hi�h煹�8�'͉ϘD:tR��Ǘ�������O�)�|:V
bO�FK�@��?i�"'��f9�=��Ck�j��u&�E{�}�����$��ϛ9��]Y1\�u!��/�h��Qk	f�#'⶜g8y#g�jP¥�O^�tP���6�L$�Ô�4pÍf�z��,�K��F��6e�5 ��1�Z����N�j3�V	jW��W�Q�>\>� ����5�w���D���4'x���A�����Ij�H�Lċ�X�K��V�!�;H�L�u1�� �M3_�\���BB��[z��N�~��