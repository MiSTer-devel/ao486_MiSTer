��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ� t���=?�t �@U�?2.r�n9@
t!`�HX��ӻ���͌�S�]8VǼ���T�T1��W��g
uNE�-w-V�_�2VM3i:�����l�s<�)Օ�>,���}M8�
-EAWL�b�Rޞi�~s�f���C����h�::� ��nd���^"���2�+��%�m��ui�hD�m޳��d��Z�s�s�˕��A���ŀ�8u��r K�0�|"�(Y��4�R�-���̞N9������5��M�����%o��`��=�*�<�B��n%�\�q� �0�cr0^�V:O�y�L���P]
nQ���<���S�O,iE4˃�n�S���a���]67��,���XU2�\�ʿ���C6޾�V�m\}�(�"3�EA`F7��u<%�k%���QPD��B�h��&O�2D��{�3|�sή�����6	bF�{dY�r��]��t�K�y>r��]�^Pa���vƏ�Q	1�����7�I86b�ca\�]���y�D���K�������S��}�c���'b����k�q(.�6����@��x�
��gs��@)ξ�����Vc�'X�����ħ_h�I6ocC�c�l�^RS�1wt��?�ʶk��L������7IZ�l˲�)��e��h������� ;�a�����C�	��gaK�Md5/�/�urT������]��Sh��ׁ�~7+���ʔ%�Y꜄�WUV8�02VP��:wn9q -���|U�Gn�b��T��*M�(�-��
\��������a��
Н�㬴 �c�L!�y��?�F�-s�������߿��W?��4��5�"����ZI� t���Z��1�'J��<�Ї���TV,m���o@���jV���$�5����0�:�3X���"o��h
�}U,���˲�)�ǘ��]�˖x�>̻�4��ĸ�ҽz�x��E2����))= �ݩ�h!���J;ڬ|@���tvD��e8��o�F���e��r}����i��2��Gq���~@�K�@���2I��t������!B)Q8����JN��pp�'FBÛ�y��H�f�����Uѣ�-���E-��������
�f7B]�23�P��p�8
֔*�:D�ЖM��`�a�O��ќS�����n8_E�n���0�?��V6N:��Ջy�i<7!-��-v��4��pS�^e����.N��?o�WZr��c��z��R3���0O��"�uIV�)�p��^�(�_���߅�������d[��܄�h�>��FU�J����w�b�����3�Vm�`՚�&�FF{��`�#F&�y� �S�XH�)���(I�ݟ}�h��I����I�,;*�%��4�r������H˷b~�X)�n�
~�ч#8a����_�iK����랓3��QC)I��e��쐾�F0�=�C�P�r	��Ӕ��-��vX^�.cqZz�X]S5v�J�Ϝ �8Ӡ��DI{�s~�f�����#I�i��S�"*�lv!��ci��R\:�EJ����F�PX˷��$
.���d�ϩ��Tm�9W��+F! �S�Ωگ��NzpYz��/���D�2L�j�o��Xn�roА�o�*.���Y��r���1�D���Ӥ<�gU��QmX,�|���� ����w��st]�b����?&�{��W�U|~BsS�V���}}�i�"�=����P@�;���wtX��Z�Z!cx��P��r���I=̟m鐎=(Ny��ކ\\b�����I�٘�q��Nܫ"'Ň��t�E�z��@�r6���Yf���ܭ� xV��\�6��'��X>����[�;�tf�����Z�s~���5D�3�x��&cnv��\\�gG��9"��1�����҉�n�㒰�ᓪ:�_�
t�G�YC}uݵ�Vѩ/����+����w�>Μ䶥xGW�+^wmꜙ�V}�yw���٪E4J1��#��@+5�[�P�����wM��}�a%���!�wP��5x��ۊ׳������a,�U�$��H���T��S�waP�+� (��� ��Cm*(2M���L��O�,���D><�DY �?Y�y�y�(� 1�Y�6ч�6�,\���ݣ�U�V/GP���� 8�d���Vc�y�l��n�GE�ռdk!J�q�6	�T�e��q�@M�~���]�����+�2E��#�]��d���8{d+tP����dwF�������Q] �r�=��|}���]"��w{Y���F�5���͌��1��@t�g��|P�<[}[�U��������&f_f�8wl�#�H�n��˳Wڟ��演o������ <i��5�2�Rkɖ{���\;l\O|�<�pn���� k@b�6!Npb��PO@�u�������1=6�Vz��=���$+g3{0�pB�aA��bS,���԰���^�V�����Ko��������n��~v�{�F�E.s	kK���F��5�/��P�����m���T�+��	�%A��k6	�0C�.�bHz�_y((t�TwG���J#U�Xׂ�o�4������\ ���P%���n��}�T͋�
���k�\sT.f{�V����>V�~p�z�a��z~J k�o=�-��������6
]p.�g[�{nVlW^�����>tK�J؁��V��2���Dlcr��������i8i;5E��x�ak�dEJ(d��X�O#�AB��t@_�i!�ʫ�GlgFӾV����E���|��?јd&Rc}���*��غ�<r�jc�d�H�r~L��\2��C�*L�=�f*$J�,E&����3��G��?ڤ%i�ў�������m����plWה�i�(9wĄ,0���~��\E��0��~�*2c(�n���R|�����q�1��Dh����G��Dt���p�iJ,�������5��~����\�r6���6�%
d6��O}j�������V��H	��*�a��[�ʵ���D��vF�%���]��ص���&�]L����~��m~��Mu�7�^���\�cL`��˺	������jI�]���z#��ݐ�g�elz#u��,��2�o��T�|�DrAg����n�A��y��أ�o��j�7�?6�_7�ǄX�kşQ�@_x�DIIǧ��x/��fR�����ϱz�FS|���ya4b�j�͝3�/���Z�'!�GVlZ}��zP��Z��˴�+�ڬٴ�dUCM���D�.����c^�+_�:𙳫���1D��/s39d-'��|�8�>.G8�籞�r[>� :���{`@V�8�����:Ө0/ʊ�qԅF�bl��X���2`E&�H.�Q�����[e�O&�k�ax�	]<I�1�>�skvsB~��>~:�ӳ���Ư�>� �����Dz<�t҅��NՓ��qU�ٿ��>�T�7���*����u�]Ҷ��u�c��"q�:m�p��P�0���g�.�%�e���/����o6�p�G�M��H[�[��]�ޓ9u
��x��-��$*���-_/�h��k��ʡ8�/��J��qccL&#������i2�Ը�J�kH?7���1�)<���Rٖ�;k{�>�����ǆ��{�^Gn��cd&�Y���߳-��t>�}�@��	v��rk���/v�zH�g�Nq�����4	`�ij��gO��C7���c(����q���fF�p�s_����9~��_��&(c���RZnc�Մ  �7��S:¤,Q��7���(��2l��`aD3��M!������5<�B�B�&�2���aM���	���g�;L<	Q�����3l���#A�����iy�0���i\�4?嵉�؃�8ލ�ݓ�Xgkr:+'�@�]ޫg ��n�+-����jf){W_N&9a,�4-��:��醵�5J�|Ȕ��:��0�ӿ4Qx��:�ׄWǳ��:�4Nk=)�vX`n��I$���m�YҮ�{]�����=(}������&RPجε�s ������z;E��ӑO���9��9<�V�C��'���N*��O+��"�qR`xT���7	Q�W	��P��%���� uu?og�FAd���#0��9�a(*K� ��N��3\�SZadG�8:�j�A�p	�܈�BlϹM(�e�PE�JMhi�|(��xT�*:X��9�T��H�n<⥁� �ia+"s1V�6F-����l[�W\��[�����9p�]A���Z7�4��#E�p��&���a9_G����A���GsA�����4ul
��2���0�:�P� ����~Ig�s>ͬ0�vy2�ϙ�+�'���yT�� ���¤U۟�t,�$tN�A͜-.��%��x�m���&?	kל<�����fk�'���x�˶X�p������F��p٥�S'��G'#$���6��wG��[�ш����yۅ�����ε��O��>�� �4���,�H����F��y�1���JЦ��,
��B���]�N��P� ��*�u�ύK�d'��v�C��m�20�vm~pj�L���NZ-6'�S�.��|�b�T)��{��6�>_<ӽ�-��g�?��*,I�J���6��hi|��W��˦V�D�Y[Gl���8]�MK3���70&���t��R��޿��:�/J?*�ܮ<�:S�}��B�D�r�4��j&=���1Xo
[�KF_V�3~���t��oRm���|�˃���RU6�r�'��� $3�mȋ�x�Nl�K˸�����օ�ߋk{���$��|n1�n� a˴�N��yZnٝ@���F1�����nxMBY-y��\*@�_��b�N�b'����!X�*�߭<	��r��鎛��3YoU�-�!m�P��R��	5AgO��DI�>j{swЎ%jUPaxQ�iR��T�H�d�1[��4y�����u�����A�/l��ߋu�e���Iw@C�c��^�UD�zP�CtaiR�Owޤ�|8�s��e8�A����q�%��.o��� ���!�% �yD�U�vu7+Pd,���a�#���}V���pKL)�����)
�!B�j�������:�% �Ƙ�u�J�7�܍� *�z�F�s�Oc_S��J�� K�o0p־�G���F���l'<�9�4��6MJ�m�0M=5r`%�o��>*�TE,<E#|������~���ω�^�*B�,B,��0X�� *A�w�5�(���&����"��2/R�)k��9jc��7�A�����+q�h^)��sB&I�5�w���ҵu�A�w�Ooٕ�ӟ?�}��|'�/~Ӕb�,� ��2�l�?lS�G(Q�p��R��b∫J�?�Hop�dґ����T�F�p�gD&�E��̊¼�E��?�nh��=��z��#�@dP�x&Nc�y M����?�
�n�[�#�q���{#˦�����������ڀ���nL\Â�=���4�˶� /sA��9A��=T4�o!�V��Ae��{S����8��N�y*2]���N��z�e���=B��7'��γ����!�h!��mKM̬�ոN��� q��I�ͭ<)�˖�`rS��GM�ʅ@�����hpݍӞҳB9>����@:��'�p:״�I�#��T��l���c��Z�q�ѫ�@�^��mPM��B��dК���gjH4$2�E��"��MN=ND��[aЗ��»��ˬ(�"nu�NR��D汨Mh�t��������m��G8 ��>K���� �7)Z�¿ԿH���L�L��\MZgہ�S�rpH����E�U"�Q�Ym��$�}��c��>��y���)������0�����̔�cA�R�����}6��6�{����Łw�]�>神��,�>�d
<`��l�]�j�};���k�v��x����Ź	�N�]*g�*<�?�R�O�!��c&a��TӰЪh�*y�~�_� �i���s%qu
�� t"��] �O�>���VF����*�I�gd�T9K�CE���c�� ͦ��v(�mk0y�xn��D#Z�8���B���
ұ�<�l!/s�;��Yw,r>�S;��콆Oǃs�Z�X���q��,�ZٸD���$�t*��.�i��&�@~Y# ��]���'�7F�n`���|��ugq�+�ȩ� �+Y�T�?��mKOU:#b{��IH���S�g��6G����Q)θ���k}Ѭ�]ӂ����`8�b;R�m��`�r�s��D?D3q6�~���jB5�)����a�������q7�C��;G7�v}�+o8��q�zA
�z"��Z��)��脲���U�֌?`7 S�KY�e�� �#�/V��󝳉O��9�d�*AeL㨼.�cg�e%l�}KE�1o!b�#�Ë�<��P�[�e����>�<)v6����.[ �j�a�4��$d��%����IP��#\O�2d�[^*_c�A�B	كR�t������[�e~ฌ�#�MV��tt��`yԞ��9^�[I�u���k��C<@e�oB2ҙ*\�#t�e��o�#��(��^t�T]��D����f�G�`X2ofb���HP���ٺ��j�o󻒓������[�;����/��i�5;~��\�,�8��ȧN�ß��H䉡������4���t��r��20u����a��r��<F�q�wC�R��d��4���5�8���G�O�ᇧ	���I-�`�ݟ�Ƿ+^}���'{��F�*$��9Q��;����\�����5�t���(��Hv|L/�Il�}���c-'[뒷��c�zl��0�y�˦.���I��C)ibwW����t�NILAH8Ä������iIn`��)S�舊i֗� q~�C��C�n�-����+¬�/�(���z�󗯅���sz��J����d�8M�.�1����I(Ԇt�gG��7�P���Yڿ�
�����7����s*�T϶ܽ�_(���{��ԛ���r�BA�܍C?�~)�.�p���j+�+�c�ö��l��@y���{��F�$�l>縶��bCO���%�r� ͞�2xnE�� N9�gM��]����U�]1q��vSvK���Wp+=E��-e�j�}!�����SIĻ.�/�`}tC���S�3����8\ ���Ƽ����+�T]=w=��=Aǅ��L��!�@�S��,��xG�*��B0rޓ�U�2q�ƍ�ʩ|��L�PU�Ǫ�6G�?�l��Lc��N�����K!��g�\+.����y=�lhaˁ����_�ߚ�%��o�� m3�;̐, ��Q�T�-Q�Π���"Sͨ�N�N�+?��G��Z�?Cu��⬛���Gj���
�v�iR�B+B���@�ˏԪ�5^=N�s�Po����5'6s�&Uɐ�P��򟏮�,�-�+�|.I��`zN��VB�1�!�QR=�xw�����/Fϧ�tOk��06V�l�ٍQk1?�>7�v�z(�;�c�]�N�!��TiyM���x�����1'*��_��3�AE�Ik�8����`CO<�� �,,"1H�^�]R{�Y��6gm�a�V����C?1S�o
$�$�w��iŰ."�}�nnz�=Ǘ>��"����r���{��/��ҜY��/�o�ZDF:���R���quzz��<�͸J�.ׇ�������P��~�z����vZ���QY.�uܽ����׺y]uj���*t�.e��aM�@�:�G��m��c�\h���ր �1џL��}7jm��΄4�&��d�@D�w�_�1]뗦�"�T+(��GmD��D�|��a�w7;X��9�$�U�gD���~ϓz���T�<5�`�}Zqp��ø��5��ʹ5�-��*"n����0%a��7���P�@��2�<��u��L�A�Rv�{³�7��)���Y!�{i�u��7�gJ��4e���\�|b�G&5ɉ}"�r��