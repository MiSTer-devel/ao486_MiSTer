��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����<	���
�^�>��}�X.�*}�1�Z����^\o�P,�b�+�s�<��8ٟd�)k%)e-�� ޳#i͌�|�*�RU��M���Uf��IH|M����{��D���vX���n�Q�׀��Ν�����$�ˉJXO���O�y|J�ڂq��' y�,�&���0sw.H�<���	���\�o8�f�[_+|m�3�\R��G�s��
��Qs_��Q��=k�1~Q��Zߋdj���Kt;�W�!W=Sb?�͹+��g��,�|;���Z�A-�$�B�1?�ز|��$�
1~Q���ע���F�E��z����2�l�"ɱS0����2�&F&�x��ćB�l��x[|I�:������E5��*m1�X.<�1�*��}l*�&A��<�I�_���Cl�D�� ��:����~���(r�T��V�)��\�uN~�G�2_�ג��KrPL����Ԍ���5g�?�qb�+�y�����{+���y�ԇ�=l�lK5�M��WTj��V0�*�Ȕ8�|{�!�֌|�Hۗo�gy3)�x�qu�iX��
�S�<������Baw�*Ɛ*q��;�������arS�^� ��mBpe�\�͚&�)���4�*	�3�W-�\d��O������곮�'���˱7=W��R|�s���V�D���'>/v�1�2	�z��F�O��%8��"?�y-HC��C�Ox5�(�YJU�V�Q��D5�^�n��m�i+)�N'@��o�G��a������t*��̺A�}�d����6�%��@�;�)��+�Q�D�A��y��|���0k5��E.Q7�ï�K� 7m��i3�x��)T>H��D`�«M�2�Y�+�S�����5b�]T�<V��Չ�͠1�bPVY-la���>.� g�K��sc�Dw����������ܸ�,y�0H�[���G�~L3`��8G&�:��X�$�ڳ8B�)\f��m���O�����ڌ�)�ɾ�r;@n{�ws	�G�C�L0�9��p�4��v���-��p����������!66{�>61G��i}�d�4P���jɎLaq1V�4�gO������xǖ��pI��nTaӤ�qU	߱��V�x�f�*e�-����[p����p��bH�Poq��o�[��D�w���j��c�%U�^�^�����;����O&���L>�;��w��|cw&�%	Ҕ�I�%��Y�p����wO�rQ�.��l�?clrT�<0�*톶�n�Q��c��FOX�U�\'uPQ&{�G��,{��d�Jr��OG��ҡ�<8��[t\z�E<9+��!l�}W�w�Ь��+�~��~r�M{���)�چ����O�V�`�c%HNQ����zl�}�s�W�;�|rr8�d_g�{��)w)��dR��,x�Z���z(����B��+�su��7�[|@<��"�ˑ��7��%;+�s��X0	8h�����&��a��դ=U�X.R�NN�V��>���w$ /v�{(NëlRYg��%(Y2�Ū4K"�������}����������9e(�"5�������BG���C(�98����M�&#]51�~�i�sb����L=@�{w�^�LM0Z[@�tK�~�F��)�o?K`��\�?��]:Y� ��.f.���ܞ��2��a�x���uO�D!�2K	��Y	�F�c�cn�������N����o(@q	��f[�>�o�r�7t3d���%,���8��w����?@Ͼ�&�$v�U� �u{`%-1`kן�Ha�;���˗_��9�;o}��N�[�g��9�����c�b8����=n*�B��!���xLk�o��wV��Ȯ����dL=�"��,ȑ��{������7Q£����b�ޅO�1��0�>���J��o>��.��ć�=�f7_lk�闍@�*��:aI�e�v�E&� �g~ɣX���~1�$DΑ�����<c*%�*e��8N�*�5�j�y�1� K~��ȶ��h�]!��k@�Y��cf#ȺP�T�dQ�����6V�NR�1Vi�2	�����F ��&�d�N��"�z�r��Ll;��9��G�ݫ#(��~�$��{'d�侻ot���fe/��#�����7-��0 ��T���y�}��<���Z)y�<a��G�Ϡ�ұ6��B�l ���Ŷ����yC_bl��۪�X�P��ZUх�F_�2z������NQ�IsyR�Oq�iw۔�<}y+<�"y�B>}q��GS�Z<��{;�|G���i}�Hlvv����E�!4�T�$�r���Z���ȫD8�n��ͥ�A�|k�]/�P9k�!O�n�������ȭ!�l}�5�(�2��t*�vw��[|�]��i��*������ʶ�:������Q9w�
6mG�v2H�Q������7����1	y�=�hc%~RJ���u[���ڃ��"6���䓁@A${�b���)u�6�S��3>��I�永b���E:h�1=��Q�l:'�l���ܚ��و^[�/v���9��fU�ܚ� bv���B���_��*���o���w�a�gз���N1��I+<ќ�(5$��qe��
�g*59ZY̊�N��K�c��q�Ύ����Y'yܟD�zfo��3ĨҲ��;�1���틌�=�de)9X0|����{�"r⏘p����k|�k
����㉘!�7���&�k�I�ٷ����E�Aޞ_�����4�����4L�8�$d7#eN9�8����q�|�Àsk�����r���T|*U�,����J�cw�qH9�樄�ʔ��G�z��Җ%Wɬ��,�f�� �%�8Z�Dy�� �s`�U�@��%����Y��a�lә!��0,y������vw#���;�;Le��mg�6\��U�ȫ��e<ݍF�ǔÎY!D:�`i~���j���Ļ?=5Ƙѻ�u��X�7���c٭�'�M��W�3zM�;xh�v�o�� ����r�+��&q7-t�~�ׁ� ������=*�E>N��)��|t1%ט++�'oE�:�2��X��T�ܦ�
m�2�>�߈�W]/,�����ZI~��5$ag��a�x�n�)�D���#�'M0������ýD(���@B<鞃��|a�|.������.�2М9Wv�����xU�Ť�(u��Kʅ���b�7�m ׌#�-����J/?�<2�6�M-d�C:�̮�,u�Yp=�
��h���Ӌ�������������]��L�t�nxo22��Mo�B����k'��嗟�� `63PJOb4z�ff�o�HU�pL?���9�pJ_����t :��	啤�-וp���J�ӳ�[�
ȧ�r��2v�p-3�*�.��v,Y�	Q> 4�8��"�`e���({ze�B����d2(=A��6l���M�I�mm� Nv)R�X\���E���A��9.����z�o�Y�G���xbc��P�A(j��c=�-Ŗ����p
|�R����n��[Ax���%�x�U��5�5T܉4���
����,�C� �qA����57r�:��`;4��n�BϹ|�|w+������#_
|
��Z:�d�i\���}���q�to��ra�ܮ#a}
�yq���C�����<d��Dr5邒>�OIK����%lR�Hc&Ù�q{-�(�Μ�Jd��}���5T��6�ю���H\>��H��\��qrfG|�K.kY�פ��3�P�?��]L�V�)�-�&Ot�P��<���F*�_!,��ծ��f�=���F������T�����.mB�I��#֤�ˇy�<J��a��)�����>&�F��{���'W�b
��as�*ɉ	��΍�! ����0J����it��J��Q0$
�x�?�/R0�T��-^��FJ���W��J�'��{��T�d�6�G�l�)f�s�\-~\�Ȳ}~���)l�X�n���{��C��O��Te�|����D��I��R�y��yv�,Kړ"��,raM�W�l(���=f��;a<i��S�kH���	��Ն�l��B�t�V�.(���V�]�dd��t;�Hn��W����h^\���Wq��%K���_3<���S�o�> ��	"
K��ކFX&(��T]��'�L�X/u�r�=:�L�Z>0��f5�&�!�3���=Mo��lD�_i�Ѳ���+����cYGC���(v�%�T�6�M"K���n�S1㿦���ri ���{H���蒥&v��G�D���"_��!�ơrT�^��%�[�����ވĩ��oP=��P����S��/�m�?ރd�F���2K��������9�ƃ.�Ċ#���*����٧=� �9u�t�8�o����5�q�KT�q
Nn.
E��P<oK��A/�L6��wx